PK   x~�X�c�-)  Ǆ    cirkitFile.json���H��_E�� �@R��}�Ru��]U(5z>H� �R�S9��u��ڗ�gZ7F*�`d��ZLg�d�����hts��?���/�r^�����v}�X-g�(��ޗ���r����-���j��{?{���N6�ߵI�n˦Z�6�2��'5�6�Ee���|⍵!�幙���^�����
$V�b���[1�T�̝�A�`�^� U0� f�*�y*f�*�y&f�*�y.f�*�y!f�*Ds� cg{ ����j�.7srUN���˚2񮫓��e�T�u�̫�Tц��Ҁ(-�$��b�("��b�("��b�("��b�("��b�("��b�("��b�("��b�u��[�D���N�D����]Dx��k�W,)�W,)�W,)�W,)�W,)�W,)�W,�Yy�KD
y�KD
y�U,) ����S,)�S,)�S,)�S,)�S,)�S,a�^;���n��,��6E��&T�Y�T�vIW�5QZWM��^0X��³���^��g/���K�����J��I��J�^~��%�}�Fr��)�=`��KΞgO�Q�x��{r/��O���n�k�N���v�s�|~��-׋������A/�lkdBk;k,۟�֐�Q��B�GKD
yE,�_yE,)�}�D��߳��B~�KD
�=L,) ���]��p�D���N������S,a�<v�%"�<v�%"�<v$��V�a�(�}�a�KǂP��vP:�ҙ����bm�#,��;���vP:���k;�����t���]��JGX�x���.��JGX:3ϰ�˰������s��r��t��3�k�k;(a���)p��Y`��ǯ���.��8� p�A��G`>~�l?p���#0���8�����_���m`�����gX>�����Y���|<l?p��#0O#��}`���`�����G`>���8�����'��~~��?,8�����G`>���8�����瘁��?�|���q`���,��x^�~���G`>���8������R���?�|��Y���4�����|<l?p���#0ϼ��`���s���C�e�~�
�8p�������|<Ol?p���#0�0��`���s����X>��~�������|\� l?p���#0WR��σ�,����~���G`>�� �8������A���?�|��`��gz��z���?<8������X���?�|��`���,���b�~���G`>�5�8�������`������|\�l?p���#0W���`���5u���X>�q5 �������|\�l?�ls�tsp���G �X>�q�(�������|Ú����8������%�}���LE_'�O�N���\)8�I�����|\��|��X��#G
N����Ӄ��8�����_��&@�S����7���N-B-k~\Hpb��꩓��}���J���� � ���ǕK'/�]4k�яK�N��W��r��8�����o8��q	�텾;XpzI~a�K�w�������N�oIzxѵ/\��_Drx'=<�/�t+�Mm/�t��Mm\�zj{�7X{mj�󷎑�(]�#�AQ��#�R��F���vF�<�sG�|���t|o�-����MnSW籁���w�%eelbٴ�C��B�6���p1���������U㝡2Z,�m�X^$yȢ3
U�u��݅s�����j~��G5?���"��*����'Ep&ic�:/�&ͅs����m]��"��(b�::v��M[dU���>�������uk��ob�I
��P��MVf��4X1�y�O}��f5�W�����GI��f2����MӃH��Ib�@B��H��%�!	�c�@B�o�"���=�$d��!	>����a�@B�a��u��H\�ƅmX�&X�F)�~�����(%ӏ���`�`�d�_,�,���L?�b��q�|��L?�b���-�~gaq���8J��C� &X��8�R2�P=�	�-,���L�H����QJ��J�aq���8J�ka��p#)��Xw�8�R�:H0&Xw�8�R�z=0&Xw�8�R�20&X��8�U��e��	ǷJE0ƕB&X��:'��s���~wm0VȄ�*��.I���[�o�\w�8�U����W^���(%�% c��q��(%��{��XG)��l�?`q��s�aL����Ǜ��x��q���1��x��q�OT�1��x
��(%�2c�����)M��s<Q��OC��
+�����]��Bb,��J*�f~<��
��+����q��*Ю����.���X@��TXc?HŮ�Ej0�`%��GQ��q��4XI��̏���U�v�`%V3?�SW�U��TX��� \hWVRa�w�u��K��th��f�*e]Ji�N�E:��d^*��C����V'�R�%Z~g^Ƕ:�
-����:����ThI���0��V'S�%Z���c[�lL��thyN��mu22Zҡ�1:����ThI�����<X���ThI���*��V'/S�%Z�s�c[�'bJ��t�2���Y��L��thy��mu�2Zҡ�|:����ThI���$��V'/S�%Z�[�c[��L��thy���mu�2Zҡ幮:����ThI����꼘����В-�=ֱ�N^�BK:�<�ZǶ:y�
-���\p�*������N^�t�2����В-��ױ�N^�BK:�\c@Ƕ:y�
-��r����e*��C�5tl����В-׮б�N^�BK:�\�CŶ^'/S�%Z�%�c[��L��th�&��mu�2Zҡ��.:����ThI��k���Vi&��T2�����e^'/S�%Z��c[��L��th����mu�2Zҡ�N:����ThI��kQ��V'/S�%Z���b۠���В-�ӱ�N^�BK:�\�LǶ:y�
-��r�6���e*��C�5�tl����В-��ӱ�R��2:yY��˂N^�BK:�\�PǶ:y�
-��rM���Li[��L��kK���0�V~~�t��#�:yY����В-��T�	�N^v�-���N^�3DLP��S�C���䪜|c�5e�]W'y�ˤ�Z�|�W��έ�<Q�Lmډ*g��NT9S�{��?}�NT	�=j�ʙ��U�ԣ���XA�xm��*gj>O�:��b��ܢ�Se0�{niթ2g��O����5G��l�x�<�T�������*C[��5��ʜYbg�L���Ճ��`���Z�Se0^|n�ũ2g��O��x���\��e�u�)�$4�J|�򤢶K����ҺjZ7�zI�R�kab���v%�Rq�.�Q*�Z��r�j��^�a�Rɮ��LnSW�3�.�wIY�G6��������r�wG�\�F�R�ڋ���1��|3��H���#�P5Y���]��(��v�r�.�T��%tyY�ќ���m���$ml^�eݤ��n�Q*W�R�u�v]�UBQD��M�����Ȫ*K���R����֭ic��*e��e��,-���\3"����򩗙oV��M�ig�>�d�/}�|��a�.o����|2��B�@B��� D !�_�"����"�����"�����"����
"���GS D !ӏ�@�@Bf;ʃ	����۰�M���R2��,,v,x���v�����(%� �0�b8��8J�l�&1L�8naq�d���&\����q��(%��0�⸅�q��َZc�`q���8J�l��1L�8naq�d�#��t�,����F�	7��J��q��(%�ec��q��(%��c��q��(%��c��q��(%�c��q��(%�Ec���aq���8J�k��`q���8J��Ø`q���8J��D����x��q����1��x��q����1�n�o��x��q��̓1��x��q���1��x
��(%�{c�����)M�G4���V�N���
+�����]S� �`%V3�OC���J*�f>��V�U��TXcޥb�A��4XI�5��T�:(��+���>��]eB �`%V3�A���J*�f>��V�U��TX�|P�
��+���;�:��NƥBK:��n��m��.��K'�"�ċt2/Zҡ�w�ul��}�В-�3�c[�L��th����da*��C�stl����В-��б�N6�BK:�<�DǶ:�
-������de*��C�s|t,��e*��C�s�tl����В-Ϲұ��1�Gb:y���ˬN^�BK:�<NǶ:y�
-���\>���e*��C�sul����В-ϭԱ�N^�BK:�<GTǶ:y�
-���\W���e*��C�svu^L���ThI�����V'/S�%Z�C�c[��L��thy.��m��VTz]Q'/s:y����ThI������V'/S�%Z�1�c[��L��th�V��mu�2Zҡ�:����ThI��kW��V'/S�%Z���b[����В-�ѱ�N^�BK:�\EǶ:y�
-��rm���e*��C�5jtl�4�Li*�N^�u�2����В-�ұ�N^�BK:�\�HǶ:y�
-��r'���e*��C˵�tl����В-��R�m���ThI��k���V'/S�%Z�q�c[��L��th�V��mu�2Zҡ�s:����ThI��k���V�ʇR���,��eA'/S�%Z�e�c[��L��th�&��mu�2Zҡ�ڒ:����ThI��kd��6���ThI��k}��V'/S�%Z�Y�c[��L����&W�����)�:�k_&M�Z�˼jMun�*gj�NT9SMv�ʙ:�U�Tޞ�r�V�D�3խ'���G=Q�L�*gj>O�:��b��ܢ�Se0�{niթ2>���T��[&t�Ƌ�-�9U�1^|n�ʩ2/>��T��[qq�Ƌϭk8�����s��dʲ�lSdIhB����IEm�tE]�uմ�z�f�
���5J���4J���4J���4J���4J��dr��:��iWu��K����8�iW���u�r�_F�\��Q*W��j�3T�L#�m�4�"�C���B�d]����(��v�r�.�T��%tyY�ќ���m���$ml^�eݤ��n�Q*W�R�u�v]�UBQD��M�����Ȫ*K���R����֭ic��*e��e��,-���\3"������&���f^�nW����m�*����X���۲n��b9_��v={�����ZN���9���[AX�������Att݋�n�Gw��;�ѭ��Vxt��n��� �'R��}F%��C�ؔ[zx'8�����ފO��;����$;��>Ah0b�L3=8��1�d@Z�r��H2���O�{r����ؕ+�ͩ^��w�������_���0�������n9��-� ����θ�'�C ��r@�NOt�1T��:�J�m�PH{�
i'C!��c(�]�?D��v�0����E��_8��A�Nx�w��X����r��^=��꺭�|��?,�٫������v-�0�H��B,a�'GB
���<	)��,�K��	��B,a�'�B
���`)���OH!�0�{�B
��پWh����h
���r�}SR����r�}WS����r�}[T����r�}_U���7�k���RD���o7^- ��5��`) �Z@x�k��[�R@x���*�0������j�U�a�obKM@xu��*��
 ��1  ��O�\/���O�\����O�\����O���S~.���!Vb��?�!=z�� ,7���uoX~�%z[�K���K�N	W[`�C,�3<�r.�	� n�r.	x� �@��kpB �# �X���� ��a��a��p �W�p �i �S���� ��O��N�OS@<jLGeP$���2$�#0��Xk�A,��b��g�bW8=���|�3�A�a��~X>��|l�Aa��b���`�*��G`�� �oPXx�X>����/Nb?,���|P������|f>(��Ӄ��G`>~]݁Fg `BB�h³x��C��:��ߩE����		M���m��H���&�w��6Dg%`BB�{�h�30!�	�r���	��Є��;چ�LHhB~wmCt�&$4!�;@T��0!�	y�چ�<LHhB�!��	��	:O��<Ţ�0!�	ybچ�<LHhB���!:O��'4�m��S���&��Xh��0!�	y"چ�<LHhB���!:O��'�_A�)`BB��C��y
��Є<qmCt�&$4!O�D��v��.t���y�C�)`BB�d[��y
��Є<QmCt�&$4!OrF����		M���6D�)`BB�A�x� Ɔ�<L���6��<LHhB�ŏ�!:O��K�m��S���&��h��0!�	��چ�(�(�<ţ���S���&�2h��0!�	��چ�<LHhB�G��!:O��k��m��S���&�:0`t�&$4!װA����		M��w�6D�)`BBr� ��y
��Є\�mCt�&$4!�lB�>k>m��t��y
��Є\+mCt�&$4�p���e+e����0����$�jx>��,f,�@��bRt&$4�p5��8}�I�I��p�F�[R���(Z ���'.9��8u�^a�A=�uY'/�y�����e��(7�n:���*��Z/�4QnPt����U��u�
Hv�r�T�A�ީR�.r6}���%��IӞXoA����R�޵��
~y!��zR�.t5U@��å��
J7O�z�p���kYv�m�,	M��<��풮�k�������_F��N\Eg��(���%w�:sM��;ѓ92F�]��F�?��	�+)�N��6uu�ͮ��y�����qdӮ�/�K��Q�/8������_�ET�w�ʘ<d���C^$y�bB�Q���K}�.�����T��?����]^i4Xaml��<)�3I�yY7ih.����οh����!�E��mR�]ݴEVUYz����_8�kZ[��Ib81�}�$�qYb(K�&+3�\L�F�����l�n��7�y�9��٘�����_�8.s���A�C��=qBF���'����L�7����7 na������[Xna����[Xn�E���t3���G![uy�l4A�D!�P�SKIf۬��o���|�s���`N6�黆���<h0Ɨ���kLB�����]�%Y<�ܷ��
>�O����l7�o�G#�"����?k�&�-:=<;������
��������$��3]�����l��l$��3=�����l��l$�pQbmO�M����c+����٤ҳ9�-#�Ѡ��l2�٘9	۳���T �NH��B2V=�+�tG�$�{7�M��f~[V�-�돘�/�]�y����'��?����G��#7��?~��Ǐ����t�Q��Q6�(�(~T<~Tp�����9�b٭淋�����4F����m�-����������o�����_��2*~�7��^ݵ�͢�s�wK���'���f�X��/��7z3���}���ۙ��\D�Y���������UW�޷���v������m�����|X�����D�h���+��ú]_��m�d�<,�+ ID���b�XE;�u9������e�d�o�1�i���K�w��4�J���-Y�|�}�����}�H7���m�e�����V�ET)�T��;�^�����|�R�2܄��t��e���b�ݛ�vo�����ao{�����h�O�{������=�c3y�ݙ��[����m{�ӽ����b���n��{�����\����b�}{^��۽�~o{�۞}��_\;b��[�6�����i��^����������n��M����·�NlQ���1�*�J�?�Ҵ�&�~�����U�����p��-YC��6i�4�m���Y�b�Gu�em(�з���sm��U	5!&zU�R�d(i�6k���v�]�=l��|7si(����ėYH��IL�Pn]�E�|{���.lY��&�>_h�3y�~q��c�&3uL�CU�hF.vrʢIlL�MaBh������z����]���r>i�3�:�I��x�.&��+k�e'T^߮��}�̶1��奈g��qf_���Eѕ�Zc�����ow�i�ǎ���ơ�8x��r�Uo7�*Y�zX����;~��K�?�a����i�����g�n���`�-n���r�(��`�u�w]t���G{de�I�tY����Ԙ윃eit�����ѥ��7]7�d)mL՞r��˚��,�Ts��6��� mC�]Ee^7g,�Ԋ�Ca�G���&yt��V]���G��`���w�_V���}�y������w�/^������{���a������}�no^lV/����_Ž�?m��nW��:���̺�k�M����/�%�޶��w���Ӎ��m������{������͛�C�X=�Lf�ҽ��1N����C�g\��~�cw�_�}������k�|Mɏy�|�:y���:�s�{��i�ӱ��<�G�.ެt3�nw�?�PX���ؼ���؏֜Ue���׫�e�z�zjs��� z��^<�]�������O��^O�1/�����}��x��\�V�͛��'U�>|ͯ���#{��E�~�]��%��~�/�KG�Qjb��pYz�g��؝��9������b������E��G��%)ue�7�5ݨ�ب�����g]�S�ޅ�������͋o���i��]p�/���c?�1S�����4�S���*l�=��%�"*���w����M�'+׽`ԓ���g}���D������|{����ۖ�郼o�����>(��I��Mܕ�������Z� ����N�����Pw�~�[�������]���7K����W��|��Wnr��Rs��e&4�Hں�Ikc����e1ڼ�Q<���.��1��"�̼߳�^���O��t��1:��x�n���`��_>���~v���\����p��vε���s��Ʌ>ﻷ�N?�����}����������B頿�����׹��ec�E�c���;��&���|�MQ���muۮ��"s��u�C��#
��ƿc���zc���K������n�����1«��H��Ç*v��^|����|���(���	7��z}��Mv�晭�b�_��K�o�m<�!i�u�gu^�r���zT?����r���O��i��/�<+ʂ�,�o��Mn,�`�4%��ã���Y?F���1�F��K��|���p��,|��?�yCq��2�,=�Aim*.<�}�.�۔���&M�z�u�猳�y�uBΤ/~X,_��~�������z�m����62_n����eH3�?f��|��e���6v��Pb���|����clc����m��_�m۱�(�6��h6�o3O߷��s���(u��Q����ݲ~�6_==��a�n6��}�����o��E����ş(/����D[�㵷||."z�r��gٜ���fe/�.}s/����}Be?�Y�/8ֻ�"ưr�����ݻ�J�}�������[������H�</����w�9��l��i���ѻ��������S��/�-�wiU��\v�П�I�!��W��u�M�����&TRE�ࠒ>�	�lLP9��l�8���ؠ����+��*'���t:\��A%���:�&��uIh7��ȹ �n᯹��`��A>��r��9�WꞱ�MO����c��ӗ6��W�����߉�M�Q�a응.|�Θ��n>N���;c׵�X��8\ȳF�]8�=�N��bԝ�p�ԝ���  �����wG4���L0+F���Y!�K:�s�>�y>�Q���E�w�	�+��b�!�*��E�<��'$����w���~f����?��w��l�^��Y?ac�^�{y_Љ�M�U�al�s>��:�ހ��ؐW��]���<Mw!t�{���1������t0��G�e�i�����L0�yiS����{���ؐ������;��l,;x|�n���e-�[0�i��t�{�@����_N��4}�^�L�LG�l�^g��
f��`�%�s\�U��3�p�3�̏��&�L�m|��u��g����&Zè���i�y���ϻ�sFv����}�����G�§֢Q��	z�z�s��ןG{�a�P�ȽNݎ>�+�۳_��Z����Z�5|+��)ܩ���yj(�Y��{�^șZ�	�:4���g�"]��Tױv���1Q��1Q�x�3�]������﻿��v�(oy��M����j���ˇ���Շo7�����O�O�PK   w~�X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   w~�X��Q"�  �  /   images/6e6351c6-f51b-4efc-b2a4-a37f35def552.png�teL�-������S�����Nq[X\�;X��ݭH�hq�"��).�/yy�n�&9s&�9N2'F]U�CA^Z�[��2ҿ��'{��P��<��(��|�����$�����r���m������wq���p��p�f�������*HKh�䜙��h˴�]�9
A�c��U�l8���]�'=�7�
0	6o�*h�9��Cw�w�nְ���<ɤ��Q��Z!�~�����R��SX0�@�ؾ@W�ܪw �X\�$�-o�>L�-UbΕ���D�K�)!�	g^T7�8RQ�P��MS�p�g�@�V���1��أ�?S�>�;e5����5��*��{b-�GQ5H�\
/"d��Ж�8�@�#��1j(���m�����#�K���B��t�>��P|�a�=
���
^�0ނ@��
�r.�!�,�F�T73�?3N�s�J�`yƿϔ�9CE�c�4XK�)}K��p�1�]hb��S��x�5�,i�6�g泏R%s�%��[ ����3�Ǹ`��i���7!ۡ�U�58·ȷ<#�"Eb�����b��cH{ְ9�2Yz�1%{�&y�v��bAMd�JG5�n�I%R�ؠ5��W���.X�� ��c�`��Jh~�+X����{�h9���^��{e��W��
�L'����p�cp����M���]�.�f���X�ږ��6�D�WA���T��봪�u��dcn�N����6Ϯi��������\)t<��4�\(t�Н���y�oEܛ��Y�D�60�!�F.�h�ʓ��g�D}�҃���ɴ��i��5���GZܘ���N�$`�Y��V�:��ŕ��ٱ�c�����:fP�u�b�σ�:Z�Ȗ�G��m�Ho��=o��6��w�7Z=�g�:�>���;�iF��;`�#� �񈅦al�w��[��W#jZ;`�M4��ߏ�OI#�:�+��O|�����b�,)�w��h���ߚ<��h�:�%wU�������Cx��Z����I���@� $�M�l�Rá�[b��j�N��3v�ף��f�D1 �X5U�k�|\��r�g�Z��������3z;��\G��M�[�)_������o��4Aw��쬪�S��� �=�3�"R���ʯ���pY� ��]g)�|��'[�,��Ħ��>\yW}=�N��P��'A�bbH��@��X��'t���+��ڢy4���F�5d9G.˨�c���o�*PB_"V{�ѐ�Y22A6�"��ߗ��l*���+��� ���v� Wj�V�,F��+;Om��+i���J��_3GR-C�$����޿�o��#V���p�Bܷ�T=~��D2f)߂v2�8��P���Z�dl&>�%�dn,�Y�5#g@�9�>��N��(�^��D��Ѕ1��p���M��YsEث���N�{=���9)ΛIϾ�y�3{��tF�X��=�I�I���uf/hr}��������3l4PO�@���i���� 5�{�����K0�|�ˇ�9a[A�=ʈ��X�oH����Q���ԫc�g��P_���3v�N g1�O��:������͵���G^�t�$��ؓT%���R���e��wE����pzu��s:\�^��V�*WQpH�E�J�e��b�?.2yéS �w� a %er�r{��I1�H����w��p�s#3�>�[�Ϡ��o<�.�C�~��n��v[���7�Β������b3�O��za�C^�T�H�,Vkf[T9r���j�	U��|Ox��!k�$J]���w�sLe�l�uk���*�=�6:bSm�~�K���*�:0�6��!+=�����8�����Όg�0dU��|d�k��c2�
���b1�߂7�"�L��\�2��UR�V��I(�8Pk]2�+���&k~tyg���b̩��������J�cm�G���$��90]���D��k!��N !6USi��7SXRm��]�٦�y��5+��W�s�u�qd��bA ڇ�s�)
�Z��Ũ�:TfP�2w'��T{�}�f�E���%R�þ�rq��4���Y��������Uj|4랻����<+t�\�>�
�B�|p�%P�%�x4r�t�%�"[��b���`�"��$1����H{VuN��C�'��J�nj��_ҳc"�O�_�tӗ�
k�ȑ�֏A�ơ�)��Ya�}RId���hj�.�+�+��w.v������[�o�"\�]xcSk�{��z]Y�$�� ���KI�6���F�+��Aݯ:���m�jR�#�1'x8�}���W��=�Sy�u���kac��c�f|¦�m�]�ˍA*��jj�.����K<8�PC�\RbOo7�7?�_�}�k�I�爰	��s���ݾ�P8��"	-�Vv�: �G�؜��T�
��nN%G#�4��5�"����\��4�D�-@sj�?��X�kz��\��1-Q���eܭCtW>X�Q���Z]P���v�X%��=��0�W�tg���=tg��~c����5��oF'�c��#dm�0su_�ŘɃeL+�'�N��5e�(MU�-���b�zW�1<A}{<��3U.FIsD�D��~B6y�ZvZV@��(��M˷�+za[P8(�fPٟ&�3PΆ�
����3Q�7�D�ȏTY۞F���w�Z�������M�� �?PXGMn/����$ئY8��o�=|oJ�5�ǘ�����`���8�7�cY��6y����ra���CR�p��
�9Y:4�e>������e�f&�)*��3���z�(�ۊ+��E�Bq�"� ��iV���iU�\�>�[K�V���I�����*�bP�+�`w]o���(ne�7�_�Uo��H0p ցa�}P�� �|v�[I8^u|x���E�x7N8����H��#K8�k\���e�	���g(w@4��S`n��
SW�~�S�/�[��C�x�f-��]��gM�4m�
_披�-����m͓�zT�˸�6.���/�Ň{�\�n����V���\��c�R�	K*������H���\�5�kӷ�=��K㓽���#M�l�����o}�`��S�|b�W���"�'�7=��W��{��]X8��d�W�׊=J�&���apT�m��֧*l�w)�ڼ�K+Ƨ2�Y��>�$iF�ZԧJ\Hp��Ū���3m�Z��Y�ڄ�t����4�+��IdH��ܕm�Ͼ��Wq}5��6Nf�#۞���
]+O?U�-�ZW�G�z2�������K��?�OЬ6��h��Q��ܭE}��>����G�
�=�;�A��V���?�'H�+�����DD1�7�ԝ�~h$�aD}�a���֮��B+0 ��8�����E��T�]�W�6������f�t��}�NZjiB��`$+��V�j��!&�o�T���n��?�?���Z�+.'$"y��0�G�W�P@$H�`G92����*S��g�m��=U�t)�?�D�������W�U�H��e�e�1͵���Az��I2�[K�EL�'��F��� �W!"�Y���X4�J@+,r�-�0��K����)d��I�O����,�ǖ5���< ��A-���G�a�#�
�F�c�]+c�=�ᒿ�|��R�y�qt"�%�>� ���_y	P�S^2��^ĆOg\,3���oKN?��a�!׺�4����|?t��!C�VRn��/�e����uk��N��XឌϞʱ��(G��w@D:�55
��$�rJ8]��N�y
�w:�P����� ��#�H�T�[�C#mި_`��1:#����/nx��o��.����e�<z�����&�`j�`�F�73cW�{�R��;�'�L�Ay�yF����﨔��CVF�4�����v'E�#d�h����[}�jlQ4��ʆ,�2el����8;GG��)��/S$D.6��}�+g^ں��iz��`c�Y�W
I�7�6�/�X��foׄ�9��R����Of�3���`�m��� !�QM��4.����N���p3E$��$��"!W��ro<����d�uh�����i�Le褾?Q%�?���:��R�q��{�E�<%>�Ňvs03�l���r=q�r3c5����`26�t�#��ы5t��K�e���{@^xIꂵ��~�<|�~�D�,neEK���A���o�Zϻ�R�����'&&����E=��������ߎ����a1e54�����{��FE`|�����<�,��m�tn_g@�v��� Ý.�ڹBN���j�B�XS`̥�}���ޱw~��*�8aG)����ʊ�����Ƙ*r��U�;�up`Y�3��Ņ0�H*(ĸ��v�����O����t��1n�pL�wvv����bD����G�X(n��[A��� �0!��h��\�<7���k��������z���^g����_wF����"M���������4v[X���h��bw�"e������H�ޯyl���J8�U��qm��؀5�4Fn�h�����L�����b4F���Q~��C�*�v�������N��{�k��A(-F@a�,�KD0E{�d�:�H.2,﷟i�0�U���7�������K7B0��{�>�ѭ��[-�����E�1�[�􈨶4���a^C��FJ2�6�}����Qutd��Ր؝W&�~�ܵ��m��d�ӡT1	w����r{4����TQe�oޯ��q�z�NW�E6x�k�&8-N�;Ϛ֞��f 0�-��h�謖�?��y�3d���|�7%�;|�s��4n�j��a3NZ��i���'��_x̀A��9d�J�yG)�%n���ȇs�B��\��e.�ز��(��"���<�k2�)D/�� 4��B����8���r�;�U��`8��#J�
�o��Fw3��겼���U������I �7��W��W��(�h�WlNEǯ��Ru����,p$վ>l<�r�6Y����%bo�ȓ�z��dK~���N�4��C��x%PlE��e���y��s(��͌wk �|�{����M���ŜK��yO��/3�fQ��MεiB��Zv5���hi�|L��ݟ�s�����o��/��ֿ�_.���fQ��R��{X�1���j�9�����.�=X8��vF/��2ҳ�;j�x<��[�g+�]GSV�C#O�f�:vP����jnn*V�D�cm9���:���z�����b�TA�jNfv��B��Ě��1��)qˡD��hd�F���~�X�b+g}�Pj-�rjۚ/U	�� ����8*�����+�`�+W�O�V�ӁOO��� !1����_�U(�۔���R|���l�t�y'�D0�IQ�;z�#>��2��3����X���-L��d�D�"ڕ�0������_��}){A��$C�7Wh����X�t�0�(x�h\���1A���x��'N�'�7ʟ��V
�6��5�țئ�yV�b��Kz�)N���t��ά0�����q�'��i�������$��ZǨ�
��^�y������Q�璤|]o>+�1��G�;�^�+�P�獿%�mc���20�I�9T��?��y��O�a �)ۚ;=��-����v���a�|M3�1�'EFh!%/�3��^�΂�*QڊF��A;���c���1��� `, D���h�V�hK5n�\������Xש��KS?��:�iҋFd)���M:>z��h[����g'��:�'�vRbup �*�n�	�TRKw� ������}sa'���A��ōy�	�	HBsg��ߴ�[~Sj�m��U��U��{�x.�4jjX���2]�U��v'�~�ц��f�ϫ)���ch%.mZ���u:e��;����[�m[V����xN ź% �G¥4�����������;h�E��Hnw�y��}���:����^����x^���)b+��WF��7̪����.2TL ����z��Z��E���+�ʋw���o�/�^�l��R!e�|��&~��祯����o�'�����i��U�z���-��:g�g\��I������A�%�0�!49�w�y���"'����!��`m��R8ņ���($�
��g�{�[7M^�Zu3k��NH�L�K���Ų+�$2�|�.tݷ�?7�}�v�ܾ�}8� wv��#��|�^���US8��l��7���X"i�Miݲ�C�U�]�S��f���?���?+�0�p"*��3�a`s��@:��w�k�1�/��?%6��S<N���M���L墴|�j����R�����LO��R�/N�:m7k�(����: +�)l�&��+�p��
�dN ��,d"�A�b�����H��;���h?���YK�da���X���z�=�j��<�g�.��yE�T�y�gk�5G?�-��X2�bTC։��)L�v�2��/�N�k�ap/��0U�#;��2�kUM%������
Qql[\l�W���?�{l��B�9m��%7��o�q�rL���À���Tl��gۥ�%�H���<Dţ�7�OG�<=ǿ\G]�xm���kRxa��&X�b/����M�9�� �@������9�x2�Ԕ��}^DR���@�A�Zb�|j���j4���W�U}޽ă1C�E��-S��=���W�����be���i��l~6�`~�,~(��Q��#}c>�����$�tU^ј(��i��
?���M_,U�"殗�����:z}}EO�0>��Ӕ�?�'�gSqyHڢ��C�ٜ�@��h�+k����K�-n�3� �c����w���\+�	c2�R��z���й�������T1q'CJFɅ�O,���#��ݓ���+����̝�0�½��+�gEr�LT��3�W^�j&IܿR�Q���4�PK   x~�X�x�LA �h /   images/7f6d2589-4c6d-4619-9f3b-04025fafdd34.png�y8��6�TJ�2TR!ɸQ���I���Y�AB�̳Ȕ"I6��P$2�6�!�y��k���������8��i���׺�5��y�uo�˚J�h�b0�}*��:��3f�N��������ʕ����6�Lc����pV��(��]���l�
�q6w�oٛa����ܳ�t0�ekv���<�(}�9�Q��p�%n�[�ů�����1_뱧�I�,�(�(v�\&��(�<�{0H�,B���Ldt`a��+<[ƺE�M�y,*0�fg�'?zw��X���)K1�M�8��Ʊ9��A�A_���&�#+qS�����,o��;�����:S}U����^ۘ���m���T.�pm�Ϊ�p��X�Q?�e�}kd��@��U���5�Q	=y,����̻�&�w1�Ff��+��w?�{��3F��K7�a������B��a?@�@�8�nD_)��-���w���[2T���h)g�ϥ�^�9<�j����#��us��R���
/���_>!�o8�.H�Kx�,;�}'G��LϢP����Zh7q=��}���8B�H��D
}b���� ��2���3��Y��T�q�3�����1�ơ�Q�Z����u�ݍa}F^���Q�dw����@�+�E�l%�&ѧ�p�����|q��h+�I�oQ$EE�'ҭ�����#���B2jTI��s{����j0�yN>�dw����9k.9

?r;@ZI��3"����>�,��-% j5ZV��>ǚB�����/�!�h���y��E���e�7��c'�,���3��jXjR�$ZJ����Gx�X�V����,�p�Y���o �婗���_9����h�l��� �#�[$k}���������R�(a��q��%�?<H�B^�sK	���@2�>jt�z��(i̚�����*�"��X,y$�k����o�w30Z�?1t3$�n?|���~$�<��,E��l�c�%i��	�Y�f�
���E���R09�0��D�#x�Sd���w1����2j)��!r\"D>�s�z��픋�EΘ
lyܤkψ'�#�=z���n�k�S4��kz��N��<���L�k�Ǒ;Բqd7q�"yV��Q/ꥍm�S5e1L��ٶ�e�=���5�MYخʳ��r�]��,Ob�k�b�$��-��y�}~�A��5��%M�4�{Z6Dv��(��)H��u�<��ٖ�n"׶�4�K�ɞ�,�n�?Z�:��1dt괌�v���M�G_ȋ�� �t�PCr��omԨ�<�����Ç����������s?r�Eز�ǜM�Hv���L^ʑ���E�j�]��;jD�߰�Y���3wmߚ$��(8�w���z;/yu��0�����+.��%��&wK�~������xX����$GcjR�����/��(����^=#�p������[J��[����E,��M��kQ\2�ߤ�F���7�~����M:������I��4��7iXA�3�/'A��3�ۏ;�������P��df3�豄�ϴ3�<b.��ot�`�.ѪV�8
V�7��l�{N�7�D�@�/���0�J�.�l��ٕ|3�����<�>Ђu�o�_}�Z�f����ׯ_-mm�-�j�99[}!چ�~��ʷ�Fg�{�����m���WrM�>�%`�M:�s-;�;��,��>�|��>dP`�{��w�����B�ysB[(��J��[XF�����^V�#�KS\p9FQ��&�B�:��|����y���3Q���QK���f��c?��z�N
E�U�>�&')899�{-���TRTSS���5����'�eu�=���TɒQ���ܻ-�׊���	�vj��8�o��fff�C/��[��.<�PE���۶<�N�/&jY�*}�~�}���.���j\�1�Xi�c�sn|ܿ��j{9�ş������/���z�\�}p
��9%�׋[�z�-���q�Wh!P8==�:Nw���ǂ%�Fedd(ci���YZ:��>g1i����z�Wvã����5��yk�yٕ8�¾�\����/`�>�%�dQ��76a��g�����-�W�Ъ)uZSvc>#+KKjN��v������\���6>u�n���e���&�qv�l��i	�.E��&D��o�\�,��H�֯��uKI
 L�WVf����D��T�hW����
�#jZ�d9Z�4��l�F~
K�h9k���2M2k��E��#��g���}�o"3��������O����t�wii'��*~�r���Kt*�,�U��eu,}P�{�)??5ᒛD����p��oQ���3�#�����ހ%Dv�E=�lMʝ���u�_+���'�11�P����6R	;4F�\#~d>u���SE#(=Ҫ�N�Ќc=}�tf:����}FvkN6����6�2/o��M �&#���<'ԣ��٫�>�1�QB�������	.�,Y9����pr5-���ۭG�k�*\��{���R���7�ɌQ�$����s�ÑƜ�q���I��)[�<8�ֻ%�H�v�[q.oِC�J?$rG�ƃ.3m�X7$�1�a�:������~W���K%��������l�@��؛P-RG����7Cph��X���~���5��%^�䣗�V��3��.rR��@�KV0	K�1	\}�p�kRϱ��aN���ɮ�'�zˍ��*<�ΐ����˃����Â%�:��C2JK��5�dҲ�ϔ�|���LO8IB���P�˃!!���Q��I5/�զX��=P��ZiA�t�jfgS�ҙ yGvՋ�W<j�lB��	7=�j,�@w�aú9z������H�.�{�X�dA/�M�����(e-��h5r�l��s.Y���-�K�*�D�maaaҖ���-G��kǉ����W4kȼy��dv��[���sH������g[I���I�/8�+�P�,j�2o>>����M�"����	�ǻ�����)� \8.�ë�T�*��*�����G�r��UH���dZ�C!�8q��*9x)wt� ��(�>h�sʽ%Ǹ�����_�n��[4	�F]���G?��c����)�q["�o�����z���oq"�Gt�_z���=z�P+�����.�ҥ�)����J^��e�z0��y��~�x���uwQ�B�1W�������}�W��tu~�S�i!�#�$=�gs�x��m~�%ْ���v��.�������Jg<��F}�WGG�su^�������:o	��>'��n�{4µ)��/-6��޸����S(l_o��L��`+h��۩����K�+z��C�tenkȜ�j��іLsR��g�r��k?C�2��L+G�u�\����4���G��jq">'Q�&�����K�-�%A����h�|������:�h�y�����,O	���_108ܻ�W����� Ɣ54���IjHB�8�y����g�j6?�Gl�=ۗU�G؉k>�c۵��|}ɍ#Y��x�v�*�M�:�.ɦ���8��\9�o�]x�GG���'��H2�d�7)$�/3����]�K���h�̗����e��l$05��`�-J8��� ���߄����^��$��AE�q6�#%���k�Jg�I�!Y��]#�xV�0��E����m"$�n�s��ߘo�5�avy���?~0ѹ}�ʱ�,�������d����c�����ǉ/�]�32i�.Fe�m~A�2V�>�8��|�Dv#�*����ں��n;הm��v�=-���8׿љ�B`ja۾r����Z_�i���<,g+Hi� ZPu��X�:j��MPU�P�咑��%�F�k��irf&��^��}FC Y7��y�و������RasjB��B �=�	`��� q[ҵ�D:�T�<ӽr�zyfpۦ٤��cgJ���rx�ϴ|q��^�4�	T�0�o�Q5�V�R��E7)�m��! ��>�LW�	�a�MT/�kRÒȬr�fm��H��������K� �đ�"M��o���An�c� �(!������UK�!_DaMQRŒjE�j�37�w����K6	��R�͍���S`3ζ�QQ�ե�0˱ o�{�	���	ؔ�����=	�	&ʁ��g�y�H&0�(**_M��/�����ʔ��t%�$�<?J���7�e7�323!� 2O�3I7k��p�L���?Ic�g�?�@�,o�����_{M�F�	�K��?�;?��Y��|1v�K���bg������ϟk�up6�>Cx����
��k�B��Dl)qw6��ܲ��i�qG����M�����)���g�:�&Qz��ף����L�N�(�yonX� ��)qw��~��� ns�RFbsyay�yv���s��
9F%�x�'A Ds6F
� y�.r�g2�;?�~/�0i7���z�K�.�� �ω�)�ym�}�H�D���)@N��٦�1���Ⱥ�pS`(\ŜP����}��	!ǹa����P�G_�H����?y�drI	v!��	<���*��9�.��)�b���I$9N�J#z��w�r�kw��LO]�4z�;�huq����Rw����t�%�K������� ~�{��c��}��
����k�r��p�:�K9o)岫���#鮅��0���}u14+���時JV��e�a 5����s��l���̧�3
\}��|���x2$, ��W��Ȝ�'=� J�, ow�a�NV4����\�b�Vȹq�����-��c�̄f���q��q��-<G.���gB��Acf�_>���ӱ���ޛ�Q"�0=��W��)QQQ��__��x��;|&!r(Ĩᢻ�;2�$hd��N�<��83''�Jm%&��5廅�������MyGC�AM		�����>>�������M7h���C�ja���!����(����5��Jz��&��;ߞA��js�	GY+�>]5��A C�e��D��;�������<��E��)<N�����[���uij�����y ��W&����}@��D�T��ϓ_l�.�Hi`^*R����-FT ܊f@t9�M���� #��P��$�������ѓ!��a�GK�65����hI���m�Г+廙>0�ք�o(�I����z�9~�l�ci�� � �}��rJW-��gg�)�'����.O�'�H�i������� ��Qæ�v������<���u���_�Jˮ���5�<r�8,n{s}�l�}�����L�4�.�{0�گVb$��[)�9�Ed��?[�d�xV�"�ϸ���
�&�����*���7	�^�����^p闧^�|��0\s�4�U��bW����Ijw����!Ӻ࠼f)Igb��k��Y���z����������B	�<,@g�S/ևxͧ��{_��̧k�2� 0��U��r���M5�ֲRH?&??����d��3��[ӵB긼���4������bg�2�x�^�G�`�d�֡馨����{�λ��g���7[�f�����
�V?7���>0�L���cU��A����i?�j����̄���#��Ny$��ҪA�����н>�+KV=ʣ�P�P���B����6��֧�]N;�Ez��q���W��v=�#5���Gg��E���Z����SQ"� �rsNv��A�7'i�"�r��:����f
�=� �%9i"�K��R�H�/���\�3%�?YE-��x�u1 ջ<���t�ئ�8����L��h79�X<��\+��������6�:�!�n��n��A�<��1]��o
&s����t�X����?�����`���=�T�p�}FI�#����o��<^��������D;e��T����h(ڦ��@�y���2l�ۿ�_�`�_w�'�����R�X�e���h{�B��N?�M�+S�����F���ma|���נ�$��iq��A�/DM:rʰ��tͺ����Hh�(���(�����!���U�C�x���&I���X�����:��ə`��ΨDr�]�2 �X1A��~\^.�ΟOC�^a� -.��~�e�NV`>���Ғ��u����{��WWW�B������A�H=rX�<�j~a��W$���2q�n�l]Ůȍ^���_������/�kyX/��{��,��q�@�_��"�х\��1;�\�Rz�6<	*�Yf�j}���64I�,��ڧ����R;�bɫ�� ��������x���,�t�8�� j�h�O�8��k��1��)cS&vw��9s�x��M�k.2��k1oy.qk�T�Yc��7���X�L�=� D�&2a`�-b���íK��?Հn-����� kQҮ��lfu�i�G��Nb ��+��z��w�~�.N�#h����B�����Ѓe���P���K����F�=G�
m:e�\p|z�������'���F�R��7yk��u(Z���q��⬅v������.�\��\f�if��/�����&��gv�k��)�����9�TQ��5a��}"XMm�`"�� ��9�o��-~�o�)�I�L�9�bx������T��=	�怽�h�����4�)a�v�om����P�(|PB@�Q'	E3�5o��G� ��A1 �ц��[Uɠj���o�̽ך�&�`�gIҌ�LM(�� :P�F(
�t��-
1]\�}���������sN�m�rM<����$-�Q�~?�`��choY�15td���jG
p�̑܈C��XWw%1�r�e�Ei�E�Kk��������K��0�cTn,��v�|��Ȧj/@���k���bA�8ڐ�{���b�@�f|�-������*�M�ҹ�)y��棻���q���3�@;�ze���2@z=���@����x�kc� h��]&�|p�rK��ּ�#�3rN��|?Э{�w}&H㺭5�-�҅�6
jjj���ㅷ��6��@	�c��t }n��ɧ�3��RMnW ��H �O�3��ڿ���Ŭw�N��Dx��RY�,�_˷��KVY�!���a��~�픽���
������̵2/O��`P. hNF���3ξ�_Ht��"�=�jM������+�e�;�o�v�����$�d2X�S�`��Cvk�yP�xE5���{�B|��sZŘ��@����F�%3�# ���"�mUbǯ/�6���j<���L��}��E������Ht!챎�!���n�S�������#��Cr3$	@<	�8`5�y9֮3�1(���Ę��?:cX��N��>q���~	���P�Vm0��@�@�3�����P
d> $
|�[E��(�Y��!9�t�O�����l�0m @Pu�1P�5���i	�P;wj!rk]��٪�[��=�������Åv��XZ_�dw_����Z�J��f�ԻN�{��3�Ro���������)F޲;��^���!�'''���J��9-[��ې���g��� ,��5�ڏw� 5������1�nά!ԙ�p�^ �� ��э���#a����NS�����e"�5�3E��m���4�!�X����z�%������..�ZEߡ��7��8��F��CٙT��6�8n�$�k<]��k5�8Xfu��ˑ��N�h���njN��o��5I	.0.>�V���y&=}��sș��V�MWw�5��/}	�@^��֥'�T�n"�|��܏ZtRX�X}���qY��mll|9QN��������\S �"��+��*�Nh�۪}䳌c��k�4{o�I��]��%CdVﶵ��ae<���E�VH�������!lM�����f�|�ʊ������n��B�ibw��ѹ�����2]�($�9��y���$"衎6��,������!���f�hG���Ͳ�n�)^�����:�:2����Abqb����_9^L�E��)��'�e|���90h�~(k|.٠�Z�V�V��r���o�e#/��"u��a�}$b�+#?_�����G��{��eh#j����Q*.Z�u_�F�[�6[��j�؋�����v��K5]y��g�!���@���*�YFf�L��	b!�[����h�ه��Z����@���L�%"���8��Swy���sn%����� ��X_�>�ۛ4�i�Z	���܇���LzBÀ��J��@���@5)#ו�(0>!_ 6L!�3�=���ՠ�Cg�
��cY��
Π��ݞq~�'}	ޏ�<��W��ʶ<�C9(��h�:��t"T���r�ֵ�;�:�����!ІigK�0.�Y���Bh/����D8�z���e��)�\1<H[D|��lY���.���|��mi���;��t�.Ҿ�b�G�Ɓw�
v��pb%��ƌ��(�Kp�vv^���P��Sz(�r�q��Sw�1=� ���R��ɵ���SK���S�[���&��*���Vt�6d`�w��Ǥ�q��3�#ho�yE�\b�n;�Hgq@Ϣ�v��Wo����V.=�럕]t�N��
+�S����_��3�q��<U�a��ʋK����b��ć*Tf���ӨIq8��Y�c}m��;*8� �}w\j��A�?�"h���
"�ouĮ���
���jP܉ӦxFq���,�A��۬��]r�.���[�v_�S�ݢvn�C{ܧ4l��&�օf&H���S��lm,��|�Br��y�+��є��������@nMחgv���:�gɆ�Hp�� O��LWPX�p��*A�C��܊h�Ym\�ȩ:`O�iS�i�H�dT��3)�'������,ҭ�������,��ؔw��(Q�&s�8�o���3�{ة�,>{&��&�<�/��Ik�^���R��)`Z����|�Á�l����6ݳ>����F���}~�O��z����L�����t�`r�������-侓i>M���ls!���>��{��dm"`:�Qt8��u.��h���ngc��jT_e+�?83;w;��b���~��ѵ��پ����x�}���	��;�It.[3g������������2���#�vC��3� ���x���'����n�6Vk"K�S�W)c���p7T�Q	%��S����!���нnx.�"exÅ,�WEEEm"���Z�ń����0�����LNkx���u����e�z���*J>Lv�r��C��a�h�Q �����<�[*�x�a�P�0�/��(�o�)r�7�R�S��N86^s�w--����Τ
zf��J�5*q�n%�醤ڙ�ۃ����.�w���,�(�RO���8���m�#8{v}���k|���ɓ{��/�c;�Q7x�GM,Y2����H#B�N�U�PS*]��ar��r� \V��s#�+%���]�we�'d,p���B~`���w[u~8��:/Iz�^?�@v�㥑���,��s���n�.�<u��AI�I�>����x��-���1��.�6?Z���']W".�ІC{�aokĜ�
�pG����7�N��,� ����� f����2�v'�; Y��/ڷځx	d��t9)Tbd���E��v�D��8S8�
�Տ�V����>���:H�G�>�cF2�^�W���A/a��w^�U�� �A�FH�0л��ҵW��s�D�)Z�Q.轞!���@t��J2L�F�=�6�l6�+w���l��\���-�����~45�(`�1�Wj+#%8 ״l"@Q2i�ag``�6�А9@#Ӈ��u�@p+>�
�G�NtC/ ���0����d' Y+,��i�5]K=J��;kOg`��t�����{5�T����o���Z���_{��-�B`#��P���!If�M���R:틎J�N�۷/��bQh)�y.g�y4aq�u��@���ɩ��3�4a*��g��\ˠ%�rb���8���ɬ���aH��x��;�c� ���qMj��Ԧ�*�ÊH��b+ �@7(��y"��*M�����'rU�45l�WJ��5�k��^�7�G郎�$&� Ϫ1�	`�.�S ����v���2�FY��+#������a�?	�x����Zu},�w�TD���I�pn��t��7Q�� 1�v�-@�d��G�<KYz����W0)����ǡK~t�ƚ7d��k�)[�F���#�kTzm"O��C��F���<:��q6�'�ywjbD-u��$��#�}������K�	����E.(-.��50���`nn��v�x�Ћ��4%�Ê��/���!���wa�#c�M�8��;E���|j_f��m�M�my�����tn\����^��~@��[ij�ZƏ3���(F�k����{���W����9��!��kR�j_+�7��(+;5|X�z[b�aOx��:Ұ�4u��7$���1�ZF�ڨ?��]j@��� 0E�p8��!��� /����#�e.�
�,]NVV�����_qc�G�K�~g����%��%jy�����7ޖ�	�GR�=<<�[��uR����י@��bSn��C_�vw��'��v�'�T���9�΅���]p�߅o�@�PP�	 �)h�e�&�=��xɭ�؜�����9ea�_����1�-��ihh��$�ͻ���j
!)�U"ؒ��$l����_bk&.i*�D�0k�C5N�z���M��U�fvH)h�`�Iˏ}Rժ�h�tu<�GMƱJ�������f6P�m����0 zu��.�L����� ��w��gh��.��7\��R 1�T�Z7�>��Z��A���	����'_�W|�Nq���"���'�)��D��$�2Z(���6z����)�O�H��xf����|�>�/�� O�}���i:|��2�!��lu>6rO��GR
6�]���_��>����ǩ�"�B(1r�G�R��zh�ˠ7��w5[��g�b1tWez&��Bo�.ɣN�i4,u(@{�H�+rw��vLOweE����|�_�% �q��=�\g�_hO�c�ǵ�t��|��Wt�		.�5�X����DO������9e	n ���;|�D5����zC�U"�����6�/�vN�T�'F;���_+�:L��e��@����e�d�QL���rYCx��� #�LX�V	�����ъ���Z�L�6E�0�~'� mGF
pƫ�7��hw�Eo��kM�{��2z��UC�e@��u���L�A^�ߖ�=x�{s*��?$������w�^ul�%qJ�j
z���+�{8���	<���֧	Ԇ|k��+5��$P<H�07Ŗٿ�MW�g�����{��t{׸�'E��qG=z�!�+ű#��$)$G|�]ai���4��E�oX�����������WQ1P�}0L������s�xҟ���qw�i�-p�⬎�@OΜ�T�[��1�v�R��~[�܃���{���X��~ĘK����%)��$0��$z���7��::"?�8/N��cݯ�^�z��{� _�E~mh�Tc��۵���~�z�-�Ru���%��G���[��D��_z__�c��ܨ���׿���2���q-((�mN��8��Wu�?~t\���*,���C�$��5#���Xi�]��o k��%o_�� .VUU=�q�(�=]�#��E��ף�D�#��ݶL��5e�������H:
�+��uH>���]�=G�<�%ͺ2k֪m�+�CJ��6l|���&S�[f�M�)��3.7x5�~:w�I��������1�.P�8�j����F���'A@_�x����V	tR���*͔p 7�q��
��`C��>���
��>XZ��.�cǎ	#	��"���Z���x|ewV���|�~պ.1�[:A�y�sw@���_S�b9s㲹y���V%������^�n�߾m��t���1�AIѪ}÷�i^H%������q�������e.���F���^���i=U�tp�_�~�IҞ���]v��@�ʕے�Ӿ�0�8a��݂���!9��?���k(Up�;������H��ifX:8���~�*��]�O+7���\ ���磂o���kbdf��gH3�[^PDA� �uo�z�c�ҵ�sP1L ��]:ƚ=��h`}����8\.�H$���x;��,�Z�a-��S@�����F"�E�e���s��'㙪��ȴ~BI���*��'�95�K�K>4,��x��XC�����ӧOK:���1.}WZ*���x\z׉�?^�1*���N�+3,�D��=cX�fs�K�}��Ol��߿O����}'===ݶ6�6צ� �`�ˊ��o��>� xIʙ8�3���ɷ���C��.-�����~�d(�p;��1��mӋm�\p��>�52��.r��k�Q��\��!F1 &����RUUU��G�Af��)��e��8�rX��8ۍ�h�*@h��f���RRR������&}�=it� �쮍��)f�*a��'�_xL�[`w��Bxf�V0L���?�w�-,,ܛ�)���9gvv��y;@Oo{C���G7��{'Y-ќ �ld��\(�� ͡����q����j�''umlr.��>��#��Sֵ�dܐz����K@��.r�F���GRLL�]������	�Ca���!(T{hK;Z[��<��!Xg��ZGh� gȿ��ǿ��C�_�~NHH(�x���'��D�i>�v*-E)d
?@1e����-��*��(���1R:�R�4;�/����*���ӓ��h�91q�y�H���Ǳ�ٕ���v�D��K8�W��Xi���ovtr�����F�Q��K��^��K�[Pv�G�	O�߿�R��u���^�~���/��uRP�c�kIjai)6؏��C:P� �c|h�7�&��6w%%?���^��5�%qȃ�/_�8R�ѷ��
�7�'�.++�����T!f����<��z`�D������F��.7�e�Ǵ�WC%��x%�� � �hw>NK�S2$���eA$U�jv�h�4ɡ���$��}��:K�\�,�>� Y��ݝ��G�l�q.��O��������^��3뾬*�����&��3�P�����D/��d�����[ƣG���	OS=nw�M���\\:�1�{��F/�K6�3��b�8O����H����͛厧ĩCT��ȵ�=f�
�l_qG\K���S���u��0�;�>y�r�jL�L1��-�I#�re��MGAO��ط��QZ�Ƀu�9��f	�Ӊ��E?'��lr�鷓�b$9��a�m����%=_|�`�q������(���4�0��ٕ�t}��/U�|q�z��GI��۠�˷�1�F�ˑM"P���gi({��x=��m��=!�3�����4�*�G����U���w�F`e=t�����i�Vn�pS�n��� &���4��XlՓ/l(z�>�C�{c!��F*`G�o���`���]���*[�bd75e���([���]e���Ue�p3�4S<�/ip&M{��3��4zw�Y�.���.yeP6U8�F���R�\�E:���x�2����^]	#tLL����#G?��'�Y��D��ol�(߽�0M�#}3�^����*�K>ƳT>Q��>޶�=�B�fR�V��3S�?
eG��p�NZe�`��|q!p�j��r66.dZ��S��Tt������;!"����`ի4�h��^�mQ���x�<W��_����_	 ��ݩVaTHO�O�堘.������V��i�E�݌DWi:�bqTTgċEIn@|�6�IV�;R"����
��%�����^U��)�Gh}/B���Z�lǖǫ��6�-��|�TJ��d�M�י��}s�./xTqD��/��������ի0+@&i�ԆUH�^t����j��}��B�WW��%�E�����zyq�z�a0�T�HHoZs@:���MU>^�s�� �f���U--1�i�[�I@ug3=&��Pi�,�`0�A[��?�d{N�:����{���\C��h$�V��ḷ�59ʺ8\��
bѿ3��*cR,,-!�<��4�yn���#��u_�ھ	�_rg�������`X��>渦8�U'�|�|���P�����2�
��!ܘ���B\WW�D�QĄ�-�����H�fW�W�����L�L�Ç���s���-��'�xk.r�6~�bllv�	���v�g���p�����yW���s�,�l��D���s���A�u����������՝Q�o���Emz�!s!G�L�������2�+���~D�����`d�8,*���30H_EE�mVp�_d H(�?-�
�
���$�O\��24��K�jǽz��K�lh��\Z�?�|8����h�~�Nǽ��/`9��M4���O�'��l��o�H��QRUQ���E����u���#9v��;�P	�3����i�������Kp'
C���E��	� 0�:�(q���8�ʲ�i���ou��_��_�H�	d��!���kv��.<��-��v}.j�Рρ��D��W+��ʳ@��nߎ;*���"{^���w=)t!�!@������e��HA�ے��PҼw�^���A11������"ۮ��X�GdW�gP��/��~�a]�V7�ŗ���y��O�Ab���4/d8م���$1	\�"�
+�� ��Ի�%M���������t��rxhh��&������0p�4SZTϯ��Ko����f�7�#_d]'WU6��c���C}7���س8BQ�t��)J���N�ڡ���U���f�OG�HP+j6Jʀ����3�3>R�N��`D��8{;�~雒;�n�'����1����{a-i�|ˎ�vv�1�:�x�5�<�d�'�L��w+� 3�YvS�������.54� ������~��{��',�M���p���J�=$�F�6�[��¶̇�v;�m6�#ed����i�R�vne�2��:V���Ç��܏�'���:/W9�#�Z��~��$�I�+=2SǥG�^n��Wnr��%������xWW��|�p2𚙛��+�^kڽ�dx��/�A�VRSS�f;MC��m�ɻ8]�����׷�#J�s�?�e�E���7ގ[��Cz�a(�O�?��t�a���6�,G9[Ku��� EXYh}��x��&!��ZX�xz����233��g��'�|�<Fr�8�=�K�8ݔ���-�=��x\"�IyF�a��$G�ެDdhY�yk�]ɝ7���˼�ct�		��e^ha��`�)��Ǌi9�4A�(�7~��f�"����MLW���I�|ax��W��� ��=o��E@0�f������ɕ��78呧�3Ы��Μ��vP���Rd�nׁ�Z���h����A����[����^�9�*W	����t��
����|�V�*z��Ǭ1"���
ǽ7B?�'ջBW��\<S�E����k�Z
�Lr:	����|VD���(-O�J�%�3��t�2�t���s�b�i�xţ������B˦?�M��7�GN�u�C�!�m<��J���}�]\�����#^ݫW�����sT-�S������TI�_>E{cTIV��!Q�c���\%�$J\��7ڜ��W]��y����Վ�l6�;�Oa�X���ʐd�2e�{� 9J�kB�m�����̠Pu���R�/�J��֣yw��~�5'���H*i*y�����tQt'�Rr�IB]��t(�+�j�i۞�Z3z�ಎN���-u�E��Z�_ 6������ ���t����w��{�z��Ug��N�z�k����]���8Z���bx��Ol��M�y�Npօ��` ��%�=�S��`����=��u�RqZ8���,'2�zd�=�V#����r*������}j`�X���cc�R�,�\��Q��c3��@����A�F��v0�mH����ߎ�}i?[[��n�g�R�N��iW���?pZ���U7��fߋ����3޾=�=J4r��^�s6�Ybh\ܻ���t`g9vز�:�dY�5��+���v��a�����_�ӽ���w�mJ�ǿk?W�3��������=h����?�n��L&���z뵼����@.p�A�Tj,!� 4Q��l�OY�Om���� ��6��Y����r3��2�ѭ��).�~������s���t�Iϟ��X+�����h-I���ã ���|�3���s9�J���3�{�tc\��g�]���q�1%�՗$�
�q.��ʳ���p�����Wx�/�*��Ȭ��S��������q0��
pnM$Ra���כ�ֵ8�|sd_���x�~𶸘��H8v�����736^s�'�7:��� >�B��6���T�����*��V����2�-	�߻��B ��1����UUUu~~aߋ:��ꘄ�<���?�ps{�+3�7)!�gu����=�e��>��s�s�w�.]�?ĩ����ӁF�
���oL���z���GL�����{ӁxC��������h,[���[�m��{��4��sN�W�ѡ����*����l��qu6���hj�~~��o��Z��h?�p�.55���e������=LR�#u[����2K�0/��O���M�}tw8��J7��b��^*ˣ�̅��-�?��p��Խq�]��oC}�0ǎ��{(rZqz\;zתuz�Ø��?u�JUH���ԿZ���*�1�3��O���@�������13,�~�����Y��U/���5�5�"�.�G^57�74���lc��o�5������M��us�NV�ݭ�@�Gw�.?|����F�2���x���|��NIII�`9t��o"�|��P�>���n�{�Ml,����U���9�j���ʅ�v`�ʡWmco���7F\7�.�|��AZV���J@]��l4$����ٝ;�#	�}}�F��/����&\b=���O�����4^�x��}���X��]M����$��7�o�����9���Kۛ���G�צ`)�k:�_�ک��E���S�U������mc����������;��+_��@�����kud�_���N�����i߈�ߥ��/��;�%<$��ky�.�Ic|���Ǔя6H��|���B�[�T�lt���h����}�v����E�H�E+�f%�1�I��_z��c)˯�e�h�^Q���JūC�nmLe���:2�'-��k����Q����+�v驋tv���z'�U�~�Ubb���I�Kh�>���p�����m�
9w_KK����'�~L�[�������r9��i����w��;���]m��;ؚ�Ѻ�{���߿1��ϖgВ�L���|TL ���TV^�.��Ƅ9h���HJOp8�3-�8�����1�@�J�� 
�;=���΄�r�7�9h��7,</N�R�maӬg3u�A�t�e�7@��~�t�w���8�s���F�Q�r��w�{�l�l %k�M�0��e?��g����aj��;���Yg�^�r�Q����ӹ^��-���Z�M?�yƧ�\��Oa�G��[�e�""��	B�����b��������\2� �ƙ���;v`�ٺ�-��˅K�.A�R.��H�"���҇�B�c��b$.�8��&���OҌWm�ݳ2>�΄�����Xj��O˜��O�U����V���##�%iOt5�K-����ٽ���ő�{��1�!<��?�	���ZR����d�R����*��nh��53�K��2���q�5준��~���K����?�2-��'g�5�J��P���#)&�
q��p����㕀�l�,9��xL�/��.���v-t�m��Lt<���Y#ve(4F�2�¶����Tm�W]=笌g[~_��r��c��x�1ү�ӕ��m�4{��$��@�UP�p$at�#�߹�~��%Z�=�ZT�}�H�;|I��I�,�;:��
�n�O�N�7(�m���k<t�~�nx$��#�R��A=��7!L������~�(����=+utt�B��ff��mLڸ��RuF�̺���m������' �4���5&n�Ab���o��z��)O�`�
Ҝ����]]�D=W�t����~�|��E0��O	���3Ӹ)�Ofgo��)}�g�PUU�6x��=��A���	�^[�\�ޚ�B��H'�OԊ4n7ޜeA�IS�уp����{�)�_�Z���f~9l|\�Y����ڍ�c���ocbuI�͸|S�Y�4'v�߉r�ۖC]����®OW�8ze63./�>�<�^Gu���J��
-��>}���/�6��n�&<��1��NA>���'���?��M�S�f���Rڰ�J�Ç��/17o,N�IG�����d�� -_~��l+�%���갨��}E�TR$�F%$�AJ����^d�A�n�F@BZ%�[i�Bbh�}��������眽�z���k��xg�4�e�Gx��n ��/�q��(:���B"*�f� ZMǍK�?�5yr�$ғ�����$k~hhpҾQ�?�:�g�i���y�흝��2�����+�Ĵ�ROs|Ʀ�K6�9>>��J�D}�m�`������o$��8�a(�п�C�����o�¸��"q��Ys�ʝc8B��@=C##9U��!�3�`NcC	�����I� ���'�l�p+��Nq��B7�xO��4�&�������_-S�u���O|��P�2&j+��y��յ[E$�D�:���^�ӈ����� W(�g�я� ��".K��\�93OOϭ߉��a&g'nu���xQ�o�#v��P��\k~��lA��H#!��Sܠ
��~"���xo�釚%��+%�Ŷc�<�͔��ֽ��d�M��9f�X4���4�yp�njD�x�$Y����ŀǰ�����Ю�n�"�dc�������=����9�T����G>�)g�����d�vQQQ�ܮ4p�_.W  �h
��t�1ţ��KHL�\��b��9�$�'��oc8��AO)�ҁ���)�穆[����j���l,{S\��D���S�;P�7�`'�_��m�E!�̈́P�@3���t*m�U<n2�}�?��:9��q�]�	����>X�k�
 2���wѽ�P�V;�,>�f��(�T���5��mLKgHѺp��!{�ܾ%�o�������߾dg�����7��lm����2�cU�����f���7�n�:���GEU��8�[,㎬F�qĴ��+M��ii����wO�	��
�,��j�wt�j���y�qt�0@�N-ez_��������9ȟ�k{	�8��ۈB.O�37&ͻ��ꪪ�op�dnm�� �3w��;���+b=D ��kCC�@�@�*����¯�


���44���wC�.�������èS�Q�?wIJ�/sҊ���Hϲ�����>�FgNt�_����`�����7��""6B)��_�)-}��Ы	�>�X.��7�+��DI)|gu��� ����ICCy��6�ֶ�wOr�Ю֭���H���H'gAN|/.��I?����<M�k!b�{����H*�N|}7ږ�� ���M�����{���%��DW�����%��'3��q6�Z
�w޻��̵�{��h�w������˹�_:fez./3Z�`(���{ύJ������_��.#�3 p����28�-px|�g�j���	�����vGW�X�i�ѓ��3���?��֎�{��A,���c�p��R�6����#k��]]C�7yմ��n�Y��dY�g�dZQ�ѡ�W]�?��t��c��QM����%��Z�s�Nګ$�(<67f]q��S|�_��Dщ����tT܁�ܡ`���ϟ=c:0{���-��	�6�׼gde��O���uWUMG'?2�ztT�����"�#�B���	�VV(��$�T����y`y�R���$C�%Web½��/��$���`3G1yK�SV�0�ο�@�������(؆�����>�Ӥை���VWS�MO��]ktY�����R@��k_[[�ʩt�JMQ���Lni���`��� ��#�c#��0�>e+���7��ó���NtW^����M���m��yKA߿������zt~~�����HK���᫊�
O��'�P�����G>|�����e��Ƿ����6%h.&1�`|�f�_k0���������i\]Yy�[��h̎D����"M�F	�<� +;���_���2��������D��\op�iR�݀�[O�hlo�5��-�?�2��G�jw��j��_=�vpX\�-��P� �
n1�-���>��xH�����~��r"8�}QQ�~��'IM&g'�9�]v�u.Ȼ�ᒕ-�-�7Ǡp����ݻ�87@��.�Z�$1+�����s�\3Z`P���8;�s=ٽh���ͺ?������
�+���|?\nn�У�W3���j���^K���E2u��$@,Ҏ��4�r32� ���nR�8n�C�x�Oi�KU��4(�B��vCul����_B�i����c���톦?,i��K�_խ3GF&���<{6AD�,Ͽ�b`VKH�+n��rm2w[��� _b�g��3�߷ ��c4��^�Gݫ@�BD�E��*煆�z@�j�F4mA}���/��!H��Z4���9$�����~ĭ�!�V7��8]�TV�0;;\M������B�o	�+��v��^�P�M`�����{j;'�?!A���ǥ{�4�`N��>i��+��z�����t��F���$xߥ��h��!�n9hKPAtl����.�R�
��m�I�AT��g��䮢B��F�~����!�_d�8:�I<�^���i���ϻS**��G79��W�߉�"ݰ���k
��!��?p&=���oo��5��g��ל��wW���F줨>��3�sPӃ����и�q���e_�%>h����M��(08��b?x� �[}y��X���'_��zH�����P�;��r��^�wP���7��f��B_��C�Er�0�����'B�?rC)��r��� ��p�'l�N���I���Z��7��Y�c�K���ݖV� �0&�`���T*�&����sQ�'v�[��VvbE�cfy�^�p ��ە&Q`/�"�@��5����fM�}
�Y��'=�4��P8��`SׂB�@�BM$��j����Lٗ��#��D0�L�}d�W�E�j�<��FC��$7.�uD�}W	!Ӷ�ԟ�+E8���1{���Ҭ�6�1Ԅ��K-?��S�H���cPj����l��a�X�-"��:�ӥ+����=�3[o��9���V���m�����T�4���Bcaыי�F�k�����w?�6Q�CK������`]�I�S��z�9��~��c쐱�dk��T�ت��V�̔y��6��'�����.�cT|�F��?���wLM���{k��7���?��Qv����G��
݆��3���ap�g̴�4F٠�<�+����F�	�>�;Z|��\�F�_	~�:���4�iE;"[ñ��ϖmo�qF�;�1�p��C���Z��B���OY��\�n�0�Y��J2�T�!g����?����F�@�!�c�	�}m1�_x��p����oN1/�~w�|�uNC;��������݅� �γ�Z����Z����7&��� �!�I$��}USy���Ң�Qj�c�ދ���SM���	/u��iD�Y2�m��-cf��2��Xg�p�ܱ	V%񂎳�vD�q�q��?������F]{O��`��BK��W6�|��Ih:�[��g���^S�d2�����S�O��5m.�s/�zp�\f2�s��9�bj;)n�"��b:�Z�.�+s�i��[銴�%����M�&
y��
'�;^���A۷y�b�x�'��^�Y�����O��0�-��yC6ǔr�ͥ��U�sp�%$hn�O�)Ŵ�WB�S����p4��zWVk��+w���+��JO�up�P��67׌���T�5<�OF*Ũ�[�0׏�3�Ъ�9�{��}��#s��#�G9`�2�-������p�|���Rél�Á@~�x�:z��&o�:˪1S�x�Ńd�����|gmT㝥�����f��k��jzG��^E=��/@�7�����0S�&�Շ)'�I�߱����ݭ���6P����[-f𕐹;J���c�2֩D�m&�[��#~Y��j��9W�+�4|�/�I�s%/w!�.Q��堶��ր��iY�(c�F���9�f�G���ô��#J�6����QI	*5=���`�O��(�$-��Y?1P�?�W������ez���S�'��آ�nyE�(����`�,_���)K��{�W�ᢿ��u��D���<R��n$Oկ?ѾG������Tg/q�XH�4fE�s�7Q�>���^kg�E�5����A��/����b��!�;���
9��}VDm�N
�J\�"=Y� (�6���,)�uK0NM���pM~��������/��I,,�u���l�Ҿ�Lq���c�,�B��[rv�ũ)���(�5��g$b���̩�t�b�f��E.��<Q9��Ͼ�/��ng�7.;O�x�G��egL��+����E@��$m��KdD����վЛ
^�����#O�P�G�R�*5�F�{��g�D��X�A��ڎݰ���w�4i�9�_�Fx[Tl���� ;52��N~�RdYk]j��Ѷ�;�?nSӽ^�kz'S�#���ғ�R��푅c�W_ʪ3��ô�T�:qi_t㞪�cc��;� h�`�#� �����?_8u�*Wk����+ �1_-�3�d?��U?n����G�;�F�E�:��	�}��9m�끜e�Ʈ�G�ԭIӿ϶6m�p)��L�����4��jLSы��7��������E\"I�c��͛^�}OR�p��_r���1��̧K�Fq-Ef��ˠJq_'��D�-�}��-jG��uӾ:w>`F2P����).��ё�#p�E�W{��NYBB��� '�xf�ގ���ċ�O��x��H*p�N5�OYH��,����������F��K��&�ߔ�L�Q��e/�\2�e���T��ε:�yt^�3�O����$[���ܳh;�l�X��������嫐,�噜6��"#���qj*_��]僟�Sc�=��ח]`NF��z4B�M���1r	�]`��}��.)�˷f>TCX�7E�	853'G������1aB(�
1���u����IB����ަ��Q�D�E�v�-]3��f����2֠�L��W�n���w"�?$6���3ai7�9����ǌd�Jme��L^Q��g)ǐ�ȸ�?z��޺���-�M��n�r��6�F �v�;���VN��2�厎��|�+bd�}}Y�����P���%[Mi���d�^�/�r�Η�u�j�3�[�B��0��NKa�N(��6<P��j��	��RNV03��g	p>���&�r�9�:�^�a���+9��EFF�ʂH�P����)�N�Wa[B������S߻<�a>��+��w�n��6��{\�Q����j��Ŷ���6�~���X/��/Ye���i�.��Ô�gr�l<�`窼�.�?�O����}ـ��W�+�R">�D�����~��Yjg�Yn����G�����K���ښ�C���^~����ɫz,��ݾ����߹Fz;��_�;dD�=�K��^4�T�=���Sq"�?�7;��6҆��<ֹ�Ή��^�����vC-��?�'���}�w�}=~��Jrfs�����L� q�!ݽ<���6j�7?��v%����ܭu��w���T<T�km۶�&Tת��;��� ��i��rʭv�۪�C�5�\�K�Q����M�r������00�;�;���y�a�֍5��Klk4�j/9�d�����L��k-գp�[����+Ft��tEx�A�@�� ����Sk��w�|�O��݃�`���V�4ou�Q��s��.ͭ���u<�G�w��o3<G��r����^KJ��e>�x�u�{�<Z�B�m�[���B�c�s�gGA��㿦N�������f@@R���Gb&:R�i�@�b9��R�w�~�[3Fe��Y��y֔�E��la��-�ae�V��z2J^��e8:�'�SP�KQ���p�8&\�ب6�ݿ/����^��J��7��|��Q|m���O�ؕ�X�2�n��l��9)��ek�:s�F�Vf����g{�����^M�	r6��?���ͅ�G�����˴<Ot��0P�2*��?pkS�7&#�mY�(��Wi���谡m��gF�J_0Q�	��&���l�_��j���Ö3ǘ����*�'5�}V�x��n[ ��$����ϴ��//���/��ܩHa��v�]����U��S��(�A9�㽋ۯQ�?b�*��mڰz~�<�v�?�S+�Mӿ�� �ӵvg�G��m��C���J<���k�[�b�(O
��#�M�b�w�,f9
�'o� _�X��»�<�2b2�1A�����Q��5#�C.��?�_��db��yiP�\�l��SO5����e���)f���Uͦ�k����|2ԙt�?�58�w�ߝUЫ�i(H�驛���jDK$��f�7���R;5���:�}�2�E"�C*#�vzS��;z�\9.�������4�ƸBL�HL����D�������A�A������H�~2.��W�����Yl�0橐��j�!��];~v�S�����<x��!�Y^� �����(]���fj_:��a�g��>(� ��U�Ӫ��$�l�b���f>(�<�P��& l�?�k��|�ԩu��)�E�PL�UƷ����F�*��^�Jvz�´"��R�R��2�C1`[��F��t>���3yk���/��UT��i�傗�|�������L���㑥��ɲ�D�ۥ�������Y��􍈥i�^7x��GcT�>��$'�+r]�qt��fT}C֋�Ș�r���:�������v=�: r����r��!�-�I>G+��#����+���� /��>��(?��n�]}���Ԩl�2)J��>�<�W���%Q� ��u�o=�%Z�!%B���,�h������>	B�F�P��pp���O�^-����?��;�� k��i��n>K�M#p����w]!áw��e�Z���LP$�Z�BC�zS��Y���\��6-�����od6^�]�-����Z���Vl�BO�բ���Y�es��e;�Ӵ���]S�n5���<��u���g��N�1���W�/+c:��P��|�a��ٰ�tC��e��	[�fY�yN��I��u����ˬ���Ɠ#��$�0~ ;|�����\TVF�T�*���j:w�0�ؑ��K;��c�������Q��,�"��ؼ�L�j�����2Q���5Al���k��yy��^~��SHn�������5L�yB�`�����d��J�b9�����k� 3ekX���ˢ˫�� �˧GtuMxn�m���0�͍m�5��T��M� ��,�S����4۝�k��
�^��Ne[�%�}��]�����х�S�j���O��L�r����w�se�=���-E�*��[��>U{8�&K.yO͝�x�R33�o�Ó�乯�Vl�:��=�ˁ\�j[1`���D�m ��-��*�MNG�Ƕ0�wNn�$��i�o��W|�W{��9�W2�zb0��i��M����`D��bf�/��ę��у�дk���w}^2~�6cx6��?|"�*��Ԅ���{x�Pgem0,�s�'��qD�d�Z�S�v�3�"�Y�~�ŇH,��[�%d:��eX��j8":|FH�+���D܇fP��eo��W���|S�����Z��8�S����Z���u��<�?f���`�;hCK�]W-ӿhP�{��^`����q/f��%����G��EL��˚o�?�����T��c�T�+��N���my�����Ց��~b��I0��8������1=0�f�����M�c�֜���V�4>��L�[.?"�V %�)/��$dʂ�����t�s��̴$��h�T�>��5Gy;�G��9�d�#��w?�5q{2��ʓT��skt.7�z��W�EU�s�cS�r��FU�I`~��1�Vf�@�g�ć��؉��ۖL��'��A.��M�-Mu%��/\���fg�y�{�_Z�Ǆ{:�.\N�\�>�v�<��2�r�������J�R�fV:��5˟S��9Kj?ܶo\�I�3�u�OPJ����G�&'e���!�����Z��[��"�c��3�%�UYo�r�:W(�ܿ����-��uhJ���&��3|��ǒut��s�_�-�n���Ӱ�q����**�<�����{8g�6V;+'y�S�2\��r��a���TX���:��'�K`��@gc@�1�̙M�J���"�U������5b1V~�B�k-y�S���mTX�g�C��U%�GK%ѫ�俗p �O�,t�R�8��t�!ť�KG[r�_�2�y�����=*�����X�|	سoig�q7����5���`���c�񒑞 HY�ѫ�OL�W����ʗ�����u����<��ȗ�`m]�I7�%��i�@Q�ɗ?��Xq۵��*ge��s,���2�w�3)O D|,�Z.s�'�S������BQX'�o��eĴZa��Yh�)|E�G�{�A���#Ӄ"K����#�3��Rͩ��V�^ln6#?c�@[�p� +��[<V?� ��j"����{qjnנ������"[}V�''��a�:e88�R�^Q\�\i[�귂ˏK�[W���Y���Ud�Eʨ��z��%A�/����yfS(��uz:�t�V>�� ������t���ش����p#�c9�,���*�,q��>����6ߛJ����Īk�%o)�C�S��¸�^bA��!�s'�w^Bi�����ID�WvW��ˌ����%���y���~���#���B�Cu�+��ߢ��Eq�,@�؄�[>1�f =x
��3bgÐ��l�����0c�1�L_ԟ"�k �a�0��|x��:d��H��	�4�v��=��Ǝ�I�V�2��M�	�:���O;�������*0�=�Wj[���B�I��wD�v��֋�x�^<ج<��X,�'��+�Bڋ�N�OM��Iw[6F+�X�X���l7v����}[�^MJX��m
���E�P���[�J�@�v��xd�����6=���	��X��<ᩴiWT��� i�MF"�;���p�R6�Q�����.�{^.��ߪ�`�U�678��܂�Z[�q]��y���#c��,��Md@X
����8-�bf������>�''�l�A�ɟ�Z�c(J�]W>��sh�)�d�4D�~q��֧7��d�K��@&�A���9̭���7C���=b�д��4���x���I[��ulFW�-a��p$��Rk����&(�����9���N�$L�ZI��䒹`��D�g׵٫Ԇp?|��Kg���C�al�B��B{v.�0������IK�&�G��Fm��2c`_t8���2ė�Qj?�v�o#P�q���兯$��p�_�q{���� H����T�_��U��S�n�E��X,�\@��QR/��,N�dJx��E�������'Ob�3@,���� ��0%�z���R�����OP�"4���e�&��gW�9@�K�<�5m����ՠ�Rژ~å�b*��΀!<���C��(靄0IC�TSO����
ӧ�-�+f�d��w�g���$m�EBA(�A�&��~D�sP��t �0D�v�E~�j�z�V�Z�����>ؠz���8�ۇ��[��E�����0�/���B���]�~.ؒ�dR�9Hԉ�P��A�q��x�"E׋:�$�wg|Լ@Y�����7V���Hg�����f���չ��V��յc���.n�����"G[�m��	��� �j`!e�X��
�V��wv���^�͕u������9�O����(���0�!���K�t�k�����L� ëD�$��a��nx�0���̱�k�Ț�o.�`n�/Ɉא�����A���4��S�١S��C��֕<t��2'��0Y^M��O�g���C	�*#�E6��D�Z��M���y�I
������ƶ���әL�}���[���juBIt;ѢJ/���ųL*�8�9* ���
Қz���n^��J���3�j��T�1t��T��,W~��b{�ۨ$�gTB��,��q�?�~8���N�D��*m�@?��oq�2o��%�){IHq�ݾo��G����H��[͍�_�dy���4o�KV�n�@�7�ӟ`C蟘�b�Y�G�+v0��؋��|v̎�<H���ڞ�[�<<�{g*�����|�B�Hk.��d�V�ڷ��y4��DB3���[9FއnW�uTβp��w��^/�L9�;�D����߳s����6c�=ެ�诎B\�����im~"��R�|%r~Q��P,�<D�K���Ŏ)�O
�w�`o��L�Zƪ֦f7ڞ%���3Ӓ�� R�.å�9�)���E��s��������^����;�:
RM8�3��͉/�xA	���u��iXN��FF�5�v��u��G�(�;�זR��>�a��M�4�}ju��ch��)�%Jz�����#�"�AV��%�F�@�mt��&o��~V�4���.��g�:
	������
77�x�㒼��	$6�"+�Çr@sh����~{�лIɤb�{�m'��޾@��$�
���Os�|���Ђ-9/Ӊ!�����E�c��5_�Է�2�>�a��Ol�z�� �u��%���kJ�v{�7�kf&Ps�Gؠ�^XN���3�������
D��]h�5��N�԰��p�r���BIYT��P��,��#��>~��NP���c�w.����u�`�f	M8�__�P��ށH �S%��1��VkK(p'@g�g��6�-��d�k�w竧�)�0I�+�<��Jil�� �h	�f�㻕1��D�ɀ�l�\���}�"�7	|� ��lH�t�i��6sY��O�t���>Uo$���3T��`��(]����j��)�6�����Xl�Fl��wΦ�y�M�w� ;�M������Y�i̶P���m3zD1[�,� ��oVN
����'��]p�L����Ѫ�h#�I�P�A��+����ʓ��P���Dt���|hhR(����]��{W�"\���m�����X�b�nȒOh�_���	��n���P�F��?ɤ��8�x��R�rF;�&N�pS�	`Ch$��s�b�#��d���u�d}#�"eY��M87���>�r���ì�R����@% [��0Ւbw{�}�32Ђ�9�*jn\�\��{�9�яBC%E6���'܎�o�}��cv�"�����L�<@�4/?�ɫ�{�0����-�u�t1�G�o��E>�05�*�6�O�*s-�wи�F��J5��u:�-w��d��=Y6hhbc1�Ҳ���@}��w@e���0���Hn�:>m|��̂������0�������75Y�\�5��I�Er�p�l�zBӼ�fC����׭K?������%�1Y_���;��̀a� �ٳ0� h��ꋪ�P'�!�['_}��J���c�y�1��Լ�	�/����B��� w�#�R;�	#l�"L�E>@6����C��Z���5����=�ֶ��ƣ��쩟(4#ă~Z��\��m�m^�;�|��Л�@h��G]�;���@E,>uq+?�W��~�`��5�(�Qo��o
�[�;US�ո��+=R��P�tr0r}[35��0��9x�@4�s7x	KG&��V�d4�-,&��9�+� i?�Fh �q�h����[7�:2R0�@�r�x��}�;v�؇}�+0O�t�2��պN���0p�B�-�"H4�M#�]8@���q���7a53�;��c ��|�!u����O$�:ޱ� ���g�U����/���Wݜ�������ca����G��m����A`#�b�Aˑ�
RYM�՘:9�XĔ6��E��m����#H�֙��6BQ
���`���l�J��k����LZAH�r �+s[���z��o��q���z�nkIL�룠`��}�W���!���T�����/��㣓x���4��2�[��;7 �ݝ�K�(�P��5���&
�� �a�y[[�T�`�cn4.î�K0k��t�ğ�'m����.���LB%���V��$m7q�;�3�PT
<^��Xp����1i[,�UD�M)�,p���Ѱ�=�.��l�N|��T��F;�'C�Øk>���\-?��W	����`�}�S�?�Ф�iÐ�PHqJ6�oﯾ��d>��۴�0�����t���z�R�̃o����Gl�ٓ4߳&�<C��xK��ay�z��XLz��T�[��8/�v��ׯč&��4Ԏ"fp��{t%����5	I�[QW]�C�g��F�+�Y����ԑ�C5J������������'g��b���Ɲ�&��|��wj e���$��I�<<��ɬ$���f\����djrP�i�YV��N@��4��ÿJ�W�<c�ż�Z��z��-�FZRx�6MH�v���S�� ��:����+*�H��|�JMr�����(n��c'"��c��~�Zq�M�zں1(�MX}�^�Y��h��ٛ�A���H�&w���b�7.����H�U�"A�o7by缿/\L����[�q?��Ȁ���'/w�B>!q!��4���@sU��#�� I��A��BԤ����QqN���g ]���c'�+���PV�%~�"m+��}�+.y�f`�N�������~L�-�P�n*|����R�*�
TLM�'N���,,M��J�u2�����qNl�O����4M�/���=�> \Fn!.!z�XО�#��9���<YKK��콍al~��� ��Hҹ��E�~��zG"��V�ސ�D�P��}w^ARN���%�.�5)���`������C6�]?�X�3�u�A}O�%�T���X�����Ҫ@*]Z^㗴��+HJx��aP4\��@t����Ϡ4�I�X,�Ǎl�C��Ψ��C���Q�:�����]xm��	�X�i�b���ؑ<��a�K��1���Q�Ψ,q�����7��Ϻ����J�깙�h$ނOpN����h�ƌ�� �ݻ� �/�:�C�;?V�����fAX6�����
h����?�<��t��t:?]����_�����3��K<�"�(��t�9 ��V4B4#�=�t��X�E����08��(I5�Z�Ih{P������9�u�c9ϳNG76����S����Jf82�V�l��ԑN(�,g1�$&�B{�Lin��(�R-
�/�ŧ٥�^�E2Js<�������ڙ��c:挋������Xk��? E�R�qN��J7��h8�`�)���ix��m��[-��
n�c���g7o
҄��%!2H���CM:�<�ǣ��<|.,`��O�蠺���K�!?Z�A�xn"���Ԥ��d�`���˰V9�m��A��1<��.�g%qA꫱9熍�Jp51ɛ���\u��� 
�f��1�f���$���"�\���47����Dc��j���S�>#�����`@�S�b� ��(�Z�\����q�nz�_��z>1�o��;�e��T}ͦr�G<��"�ᙲ���3�砏�X�:�/���;}�8̅��φ"f4"9}$�q��n�}&!�<'�k��D�ᷳ�ux.�rl��c���t����tB)<�og~�� ]w=��Ӭm�Tch�6)��(���^̚�����Y �-�+��@Eݡ�om�ht�u �T�g�	~�R�p�ս�b� �csP������3r�N�����k*�O����pVE��w�\$@��!�4��>瀆�v���Ɠz�}����!�b¹� M
�=={Vu|�	FSQzRJXb�y��h�{.�u�[D߸U��+�Iҫ��gr]��_��inC���)F�XYg��lz�JZ�_ް�1n�ZIVoAi�1��
����)��j�F3 iO��d�i}r�"�����x�ҍ=S�#�Y��P4�vbR�X6�.�}Yt�^�Y%�A7'u���5��A_�K6#<�Ԭ5h�;��/z��C��Lik1<Aۓ������JM|����(W���̊F>LV*�����ܦ�<�S������?%�a4�w��,P��i<{�so���o�F�m��!
��&w���t��f���r�E��]�3��U8/�P��(�˫����-M�,�W�j` h�)@�M��:�'1G���W �H}�&��@^�	���Y��H��m����Ԥ0���<��AKf�Ɓ�S�-7�CZ0��\ҍ:L#��Uk0�[�r�&d��И��w�^k(���v�n��������(�()m�L�H�E�?*p��Mwfa|��C��q���܈�ޏ���E��~os�c];XұJ�w�K���n��Ex�!��0-�FW�y���o<k�!}����x�8|��a�C���^���/!���<:�����q��B��~�pt�?���}�!$��?�v5�&��E�ek����<����1{��-�S�:4��DX�'�g����/���d��ٜ~ÜZ�7z1@X"�?Q�qʧ��	(QS�g��9�EQ��i'>jM��8�L���d�piFa��B��=X��ۛ��,*4�}�,G#��g����MK��MS�������V��~�y��kS�-�񸯈�J��~�n[�:U��8|x��e�� )��"L�"�Tnr�66H��*ARʨ�/��AT�$biJ������m��2��O����k"��\o]��j��Vwr�֢�yʱmsQ�;��]	��"�B�"��"1mj� ��OF"��G�&��)�%��Sk����*ӝ_��[b�t�'5]�c>�"�r���d�plioYXĐ�)�FF�)o��`om-n�Z�6�Y���X����C���Ķ�ۿtB��lW�����U�BS�7{�=�-�C �}pn�4��`�v�J#c�Q��2��D��:m`��+W�ÄW�l���$9LO�aa� �>v6�8��CP�U[_��J����n�2)6�1UG�� �>]�E,�D?x�#��M�_q�l�!2ǆ˄�{o�"�����y��*�ԃ �32��B���N�v��Yɠ4��5T����15��<��^���: X��5�͛{L��w���ꪼ<�c>:����l^̽�vr�rC��j0Ȅr�
ٿ<�� �ص�0��8��io�X��iD/K����t{x������pSxVԼR�d޶�/�ƱG�5(��0����,Ft��|�I���U�M�B.*|����PN�����~.��#�6��Ғ́�=m���QC�������k���%ѵ��M�6�nO�
�7��B�/Ѓ�W�">��`4�[6���f�_�l��������S��]��3p>�9�@�
�J�_�M�&--@�솳��,4��1B}�p~-��[�ܣ=�r�]%O5`ߴ?�(ҸI��/�{;�X�?s7�mǂ,�@d���G�Ð�.����\Ʈ��ً^(���J�����5��	~�[�:Y���;�X˾>�2�:�j&����'��������:�����&�B(c�]z'��1����`'�U/O�LE2��ɔ �Ed��<�����n����8�/qr��;㋋�Gꇸާk��ݮ'$>�q��������B���\���P�*۱<���4;p�̝��w0{6��;c��)5>mhR��3��\-��e*�Hz ����]��IC�т��� P�gg�BTe?� ڹT� JS#��pr�����ӓ��3\�� �45�ۗ����i�$,���CQ˛�9Ғ�ŕs�~��Q���IK����������j����Ԫ�� I��`�J�G(	e�_e��j5��/�z��p��/$9����i��$�k\)U?�=+e�K/
� ��&�i�������0��F}p�>�'_��j��:PА��U^����eq<�c�R����F���i�O�d�P�@�lV�l����z�Q���Xztk�2���Xъ�b�z�_�]lJ�K��33�K}�܂��P�KĐD����R�)��%񣼟+XY޾-�ƻ��<7g��y��t��q��+C��}Y��g\D|J��
6��V�f>�L��I~V�_vFyg[����	�B���G��v<����@=����$a��N�y�{Q/��%�����R��=Bx�@���l�Sy�,����
0�P�!}4���W0�{ը�z�*3�w�{/Hl�A��O�S A���&��P�(�������C>r�CK�+i� 0r�6hh�G�B9��SW�|��Ǎo��22���t�z1M����c���
����o� ���qM��CGA��E���鳭��z�	&�T�D��o߬��vt\/�&jA��go���F&��myIg �)?��;Z뎽,=�e���w�g��=�}�A�f���+���_����L��������O#��b�n�m���g���tJ9���P�4f���b��~F�'@3Μ��ʏ�@���)k�OT���#��͍K�Ͼ�L�EA�rﻱ�<�{n�6�xl��o�X�^7
�����+���]$��|-[�V�G�����ջEW�Ȇ��^;�� t}m���7!�d0��O�::�167�Z�ns�����J�W|=g����ul�t�WL�]4NX���!V�Y����h�<��ш.�]��*)�}�v}�Zu��9e��_T��#gf�'�?�ͭ^�;��K�W*y�*p~x�p<��x@�Gm/A��US�3�~=�w�{%��$��ܙ#��}wW��������9�O��߈%�O,�}2o2��G���Uճԛ���E�G�G�/AM��nX=\��w�g��N�o�C� ���ݢ^���?�k�����	��t�'ɦ)3���yA<�������p�#<|U�sa��/#��P�SP�w�/@����6�A�Cx.����u	��r�X��N0�~H I3�M�v�Tw`WA�����-r!��?��s����:���~�X��R8S�Y#W"L?�l�%��Mn���_�,Vc+i(W�ٱ=?��ˢBu{ ����������nm����$9�[� �%p�6h���K����(�vsp����A���@�U�Ϛ�_}V4�M�W���������8�&�{�¦�E\�n�F�����Q��y� ��q��UFk)&�$L��ak#&�������T����>aEE�$|���C"3d
T��ǲk:���فi�~�����f�G,c�J3�gn�{�I�<���Ŀ��鿄��ȱtx�o���yX���_i���
x5�;!i\k���'ʸ-�T��I���%�l�Г'�g�S�A��0��|�; g�|��߉�`gp�B��+ɨjBȿ��޾e}�����G!�>� s�[!������.�o��R}k�x8}jx���o�h���W��ݿ���J��6#6���j��������wRg������&dhKFFc ��/3�Ů�;�.����4�k���4v�g�@��M�CՌ������͋��c�����FL8 iJ+)��tI7
ҝ�QDE��[�RA��@���΁��p��}�Ͻ�Z�]�����0!0?B�Peo4���-!�fM>0%,�~�����VpI����}JJ�V��$�&'ӯ��x Ƨ�"}A#�
��wT���?ߟ7NC��3w�������ބ�����*{�΀8�J^T�>��Hb��U	�W�
g9�.5c��~�e�߲��k�=�0�� �W�v,&9�j��i�>ǵ����|?��ff���ĝ�b�<���O����>�B���i��HTz\~�b�}󂥕q���?�dC{��I���Q�zI���veHR��#���YRH&�]�Aw��y�^�lW�_z��~u����UQ�i�$�P�]ii�bEa7�O 䥿�IC�`���Ҧ������~@��$&;J�Z��L�u���}9.A3?�r5��:���p:��p�t��]t������|�)2�f|Mq�;��K�]>݄�Y�iw�^�[���q��]I��Mu��h�3�p�lb���m<�5KY!Zz*�$%Ŭ�*v���QS�Eq]i=qp�4�Wڭ���ua�.M��Mk�2j�Yo��4(ޥK��x'�<�X�K���~��iKp�����I/0�6K���E	)�8Qe��7��P�V��I`��i�~-�a�~��P���"��T���MC��{��wM`�Pn�>�xw2���m��-I����z�=�e��[Vʅe�h���?�D7�ٻ5��g-+H�/�ؒ��t�{v��߿@p��Ճ������V����:���6+>{��H������ a�"I@Ӱ���"!G�S9fM㟿�H�6��1�p�]v�5���/�E���F]W5:�b�^��9�x�����o$�F\a=úͣ�4�t��m�;����;��W}��E���x/%,l9�;?���D�U��M�+���������[��{.VKm�"�9�E�Ӥ�d��9�(7��|�>ƛ�y i�X�EK�4q��2,�!1��s�1����#@��&
Ī�EZ�׎�����%`?��� ��%x�'��+�,7���ٮ�x�?��̓6ᣖj-&�G�;^��g>����bu�YL�2�p=���`�4�����;kܓOr����o`�V+ԍA�+t �[|��ȽnK�nD�N,!���I�'u:C2O�z�%�9xN�M>�\@ ���B�ՠ\A����ѕN����5P��w%��25+���m6�ל����|[�/� / 1�A�
��ptD@Ԡ%XH�6������+m�[���`�&$�P_X�k6y��jf:��ʳ����mN�}�i�cjr�2G�D"Uj-�9̞��U緿��2���$��`F{1ǋW���]�Et�__��K\�!�v��H���y��_���|�ve E�I-���I���S��$�t�����*� ��9�٤k��vBw%���k�^b���Ps���H��ډ�}*狠O/�+rWT�}��N�8
��V4��[��4HA!c�2��*S���i��J����i%��e�cY�O��g�Ҁ�9��S�n��y��t�9DZ�I�}fe����X�Ⱦe���#��~U�{�W|����Z�����ֶ�|ְ�|`it�
�.�����R��v�&�e�#�$��mN��0�/�no^���,���>��@�*�j"pl9Ѡ��O���������<��QG�㊴���0���������<�6`/1prb�f��ƗĬ��}��R�ؕ�soٵ�v�}�����Z��N��eG�܍�P묠��-y�Lc���Z�1��rs�R������D濸e0[������hiS��]�h��y�}^D������eKP/�
ar1L� ˋq�J�g���B�7'o���G��dH�6�b��7M������yy�� f8�vt��Ks�/gۿ��"��W	vo���»��:ζ�H�BDн�ZZ4��06�@t�a����z6�&���&¨�J� +��y����.�x�ɿ���k�,��6�55��g��Ũ�\���-�����M_�TW�].�i�_`��C���
�i�^��Y�Lq�W��q�l�/�3�ml������j0z�ژ3R�Lv��A�-4��C��1�d�b�!˸�n���ws;���4m��$`�"Ȩ�Έ"�;�����(�΁�
�-	��������W�윪L_q�Ǥ�p��7.�E3����f��UT�/A�Z^#��~=4��S���<��Tn{J�eg�1����_��sqQ����{]{����
���[������&�8$�x\�n�[w!7�եS}��ƾ2�f��Ru��ev��,qU����GW8��G'��׋���u�*�A$��y�<�k�}�[I�_;.5�sB[l����C m�s�g3«���ZrҴ;�5('���K�~�y-�ۯ��t��:�8
�j�0jA<�s��������v�A�*@?��M/\������Y��/2���q��3y��Qr'7�ǿ[>��5K��.2�����6X@X��@ �Y �z8���b��Wگ�.�![Q�I�$�
��J&�R%����8�������ƭH�	�� ���!��uV��0v���b����E����n���ۮuY�]ﴬj��q7�ܶ�t��W�����wd�F@PXg�+E;(Ih���ƛ&18�J�w�Z���
/�SR4�p�x.C��##T�WqT\�d���7OHHh��jjj#��$l*Ib6֔Z:�m秎��bv�ܲ2�vp]FF�u�C��b�F)DU��O�}�I��������?�#�/I��c��e]���S��"�q�����37Yb�V���A�yHU��G�-]>6�.N{7�xd�To�$����[�(�/�A�uѲ��jo"�cH>�?�uN���dzW
&\:� `]UT<Ҵ�k��������챗',���n�T�2��u��bj��W�z�A��J�04S�@�b�s=�@�k�(Z9��2�{WV�T��%=�=�Zv-�R�q4V��g���Ѩ����w���ٷ����-�+����M����sUv��QK�JjxC�@����ȯ�D�疗E�������ID�ڽߑ�#��GB����.0� �/?�]ܒf4i	9���8��[��49��3*.Es�j��W��v7���Y�D;N���M�V�0���-�z$�# �:��&�ĸ���5A�DP�0�w��AcK-�{A�H:LB?���ی�'�{��?W�<�b��=S�z�Tﾱ*�adF���
`��C�d�	��;��Y�����[�����D.~=X��*5����w���}І
��uH`yg��(IXt�m�~���RSEbHR�^lt���p�Z����n<'Uk[-{s����	�m2�[�շM��*�M/�7 �_�(v�X�ǣ��^�J����x�V�1:����F�rC�JΟaf�����{�2�������t�����_�eLͲ�_QԸons��7i��g8����;�u����.�|���.�%�F����^��׉�����9�7k`P��3�e`ז���w�rb��@��i,A�O��J����U�����~7�%�j�L7���C���S~�\:�=q�~)�x�R57���W�}^�3�$�^Lx(��BH�}�\��O=7y"��X<� ޵��g��m�.B��{n�X�/�]gF--{<��T���`i^�4��J;)A��m�j��O����(�k#���G��/ ��gBf2��+��{�K��*���P.://��K�D�<(%���a�?F��H�H�����8�nEI�ѽ{��m���m"h�#b�>������Xn�ue洄c2���Ww_"5yzne�eF��_Z��-�|��'u�����X
���1J�?b���BD��n-��Krqt���/�Y&�Û�3i��Is�#� �/shX��m�Z]m�7=A�w�?|�w�Ҏ���jz���c7�ک��c�6�� ��X���Kp�\(~��W��*8��f�/�f��/�����siX��/M�%o��u������?ߤ'Җc���|�E��^ō �T�Pʄ�YV�~����]]�%d��X�����n�~����P:�wo}$_7�%��J3�����m�[� ��J����Lt���.E0`u9����PB�������
V���N��Ŀ���7�[�*@l��w����k↋��}�D�)������Ba!�W	�o��k���[.�Dno�8�ƿ�1���N=�8��T��|؞��:��6�-�>_�	�~R���	Rh�~�\|o	�[���U1pI� f>�#�M����⨎C�����X�(S<tݞ�_�=��K)�r���H~��9y�*���J�N�r<8�Π������n1	Ά%1\Q>wN��!LE��E�~W'󭕔kW����@����t\�ѡt�!c6�E�4� q����3��VG���^��n�?�;I�iS�����^���Aaʩ�����l��������uzʳr�?�X�h���ަf,��SJ��(rv���7�-u�N���ѹ��ԭ��p�G_G,�S�%RGunk�㔔b���gս ����/WKR�r���Kz�1�쑣ʬ�&��wO�1����		��CD��K�E�L�bl���M�=�7�DT�^�U��>��;Xł�.<E��I/(KOO:{�p�ʘ,43��U^b�9�v�FP���P$�����P�*W�ʹ�q���b(Vjʞ�u,�r���m;Ոs���H2bt�+�Ù���OJ�ϼ�Z>�ZI�J��o��J��de+,�:�,��(�{��9�)H���2+�V}��C�2������g{~���͛[�"bt����h	a����Gn�^��Gos���(FF�AS�g�;o;��sP���G.���k�n���՘�py��zl�㴴Y:�������1�x��kFL�ꀛ{s�S��#6�S�<����bf�pxxUָ�A�Sd�.n�wc�qg�8߽�����3�CrncU��	{wM��
�m<��H��x�Nv9Fa�zک_�UIWW5\v{��pQ%O"���X�����9�^EX,(W0\�$�y���!�r�#�]L��u�6jpO��0��dʞ��5�"�3#��܊<4�{\O���m~�G����s-���\�@q�V�)&�y��yEZs�?i<�G�P��;M�uoC�92�`!��AW��e2@��C���cm�;?߹j]4>
�
�&�n��nz1�$��RW����U{8J��,���7I=�`����:��Ԛ�Ľ�l�/^�A�T��5��B%`�
:3�nZ_߳*qӱ�ъ���z��d���Kanp��'2t�A�6<U&��`��sK��RH���,�t3q���>5��i�l,F9�<�"�O���8����X�s{ҥ��~���S�����0����D{	�{�W �+�Դ�A��td���$������T+Х���gM	��Mm����^q\��KI'������]��xI,u�4�om0[�si�q���Ⱥ��*���"}��^�����.-�^�ty�S�&��=%��H8/]�!����͒ ����_C�F��sj�����K���m�����]�ڕ��+�2	e\�9�˶�:z�<��W̥qĊ|��4@�(Q	y:G����o$,���ѵ:U���5��`��}��XS��^Z`�omy}qt�(-縟 &���C��c������_���B�E:Ϸ�mv�x�r)�����<���l��; �?�D^~3a���nn��1���(��S 7�·�*���"�K���H��1"����� H<��0s�D����eJ��Va2�`��|���3sd
��ɓ)��ֶ/ �"�e��)�Xu3����*����h���G��ڴ.�T�I[���n�v��.	������V�ο��%[��~�aMG��E��޹�.��zV���<�z�y����p�%���1�NE('�dx��RhS��#Q宬�9��<���v��J��g�I�b�0
�)��aGe=&�G�����x�w�)'��K��An�m�-�r\���k�N�E�%�A\�';[a�}���@��b,F|ǿ����~�BB��+X���x��~@,�ۅ���zz��Nf�ҿٯ/�zwUج����AiU]��V���,����p��u~�.٢��q���k0��u@ff��F5,�������t#���*���`�0y��9I��8�B��#��#�]���~i��߰Is�]���J�����[�zX���43��-�p~�s�&d��MX$0��k�*h��)6���`�vd��(��`�����E�䂏��=�ye.���$�2�;w!H�geQ��9m�g��g�ԍMխ+�\%�S��SP���%���vLkv���Qε:�	�l��wZ���6��j��eBI*��b)
 ��+cR��L��r�3��ꁟ��m�����h�Xk��C`�i�V}�u��S�l��V� *�5۵5�G�\���5��mDP| h���K�J��W�''k^� �]�_^	�i���%c������.�LCt��-Cn�PA������ʎ>�	B��rk����O�F��u۵�����]D�1[Lx�F}�V��c4D	@7�a�G����d�T}���n��,@��$�H(~���J��\R}�>�?8Y���m��'
S^p�=����W��`�ϔ�X_�o�4.%E+{|W�-O6�z��� ���;nD�J'�������g����K��6W�OH8 Ӏ��ޟ���.����~T*��7��۳���� s�����9|=6�3�ۨ����i'|~��T�����yP9�ɨ���#�:އ���U�@^=�;�̩��dJ;$$�2O��̫��
Z�w���o� DXh4��Kߐwk?������V�����m��I�X�Ƕ�n�â� �$��E�_	�(i;Y�0���"]x���aR���|���,��jf���Щ v����h��#_��;��S�����L&�����p&eɞ�c�fAu��i����u{
�)M�ڦ%��W�tH���eE�=@��BR��� m3<��5s�*K5���d}o��5H��	����VTL\�H�U0m�g�ի�����Tl��5���}�!�5�$�o�F��9��J)�QWپ^��M[J��34Bf�ޞ�PѺ�4=��WWh������i��ǚ.ZQ�A[=�
�$��媓�[�z��W�	o����\b�<(���Ƶ�$J;눮z�?����F�x$���皎����L�bj��5<�t�,���C��e�;�o���a��J�+� ����-�*�����
�zQJqv
+���,�	�Y#���M2�S�k��_zmN��;!����:�a�a9\fo�W����g�vc��:ݖ�`�V!���k�\�;BB#u��%+�^���p��*-�/ɳ�m_Bw[,~�M�����?�����
g�@�s�����X��
-���ډ�m�Nh�Wy���9�~pMo���e����Q)q�uJ2d�G<���܇��|ƪ�gzԦ�����IKV1�QN*p.�v|䫲�_���e%�@�<�D�;�F0�Vj��7��qt+�g� ]�So��~�����9�MT������x���z��wZ1�IN�{�m���^��i#zv�C�ʬ�U��E���1YM�>��t�J�Sԙ�$��Ӿ3��- y�w�v&�<�uaI���NMȪ_�3}����&ȁ�C-����lE��O�-�������'"T!Ʉ5�=�v�.���%z�^�6��S,m/Zζ}Z��b����j{$��I|���-w�S\�����˔{r�$��{�>|�����晉�i%�;e��x_)��$$�;,L�g��b
���㸦�_N#!>��&h۪nWT���M17���PQW�/�>Ϊk"^u�j�6�l��t���/*�㊧#�&2}~gž�RD;[��dY��\�n|������nC,{qr�I}U
1$�j������"#���*ׁ���������ζ�	a�����p�[�q�O�L�1������2�m�J@$ǡҦ���N,�6�aVJY��ج�� FP�wO9�p���'�wD�}�pI�0+�����خ^zܕ:����g�."��Ţ���?R���Ր5�����jjΎnF��3		��@�o�Jj�2g��:F�l�T��������zC�Rt� F}-/���&�~��T� �T�]�v���o�c��u�� sv���1{��?c���l��a%e��S�@�0_Yž�M�E�9��lE�nB�AǬ=��F�{/Ӕ��m6v�y�OR��ǋ�R`��YC
�WQ%�?��ϐ5��ς2 �>�#s���M��8��,}{'�TQ��w�'�.����C�WAVs��z��j���z��vG��g|���Q2�
��F��$Ί��}>�RV��}�8��� �4xa������L�C��认��Q6z!��6D��@�b��Ő��0E�roO ��Ƶ��U\'~��-��� �q�[*+?/��SF��ODL�:o^E���vE&Ty�]P����{66�"��Ļ�� Q�nS��cf&
��v�pr��θV�2���칱��Y�����ܧ�7����Ą�O�B逑E&�
T��&$l��6� ���š?��V�8|��U��Q�4SN�˜3wp�VI��^+�<v�-�3��tO:�ϟ��-���$t�s��d��1� �Ò���n�zw����O�?Ǯ+�����9�^�E�EP�bB��%.���#�f�L�miF���	���v*����*N���Mհ�7�!��2���%G��̄��4��7ɓ�s������\`~Ό�#-���of�^2�{�ӳ�^�Π�愼�r��ʹa�/8[��rҲ�O�^��J?Q�6~��Bb�Zm''I���j+0���뜀����wZ6<I��g�c�D��O����4go���Bj3�۠��Ŏ9�|�9����������Y2��Tq!��x����y�Pnj���>{�?fi7c�� A�w7���5c��ɢԎ>�W�W���Ԉ��I�s1�� �Y�Ltr��s���ޟ��w۟���D0����tl��WP�L(qna#JQ�[T����X����QT��K�����32���8ﴡ�ͮ�џM�����ř�\��	��W� �^	�%��d��vM��.�3�ꎜ�������Ɠce��S�- ��ĸ⺝c3�\8���ٞ�0�=p�)D��}7^�5Ǫ�=�'9�,�r���cN2Sc�㏏�c��f�Y�94t��I��#�"Ub��(�ׂ'y���#�����v�l,2�uoo�	��VMQ��d�:���^q�}�r��a�߆,�l'LT�*���Y����v�@O�8i9��B�^Y29T/C�'��C�>����V"Q�H'\_S�6)��|6�'����V�lx� U�j�?N�=����@�t�ru"L�^��8M��C���i�Y�W�����{�i�h�|W��b��|�2uP��Τ��ukba�9�Dp7� !��9�n�+��ǻ�y(����~��a 0�� �?
�[�^v��(U�,D�ǗW�w^*-�ث!�x�L���㌯��v��<Lr���Qn(���[>2���߱:��@j4��-�؟ʅ�t�*�R�����t�l��HV��"�x�_<���(��,��j�5�Y������	6>C�*�p��{c&�XVF\��h9u���f=ty(<�_��S�4���3N
e��_�G����y���]����%&�`s8��V��������lZ����΢K�.)%%YR���2�W��k�����k�'U�~�K}�/��	 ]8�s�ū�\�#�\Q9�15LE��%�غ�����hqn��n1�����,F���m3b�&arͫp+�����1�E��`EU��ݡwWmoA�w�E(���i�1���!݂ݰk����߃g��5�U���o��kʆ�5F���rm[�̈́����`�DS�8�`a�'Ƹ��W��U\SW�4�Z�K�=�m�gi��� �c¸i�7=��.,!_@ͫ�n�}����hs]{�UF����C�~~K����ː���-J��E/jy�;�_���j���F�S�Ry49�'�k��^�/iY��ٵ��?&K޼���� ����H��?/�qʈ�['��k��ɴIo�2w���0)����4��-���㵼5���G��:)�_���ir�v�9y�	?.Т�����ɺb�:^k?Ԁ]#�n�&���_U�bcPi@�DD%b�1�m{����'��5 f fL��^@n�g�P�rWM�e���M�M�^ɒgQ�烠{w�̻��y���ˁ��OK����rHx��V�O+o)9y&���-[�O�r�� �q�m@�y�:X����d4��WVm�:&�_�y�:�X�B��'��7����3�i;8��T�I�|($�f8txa(G;4�}E�'by���~������rVm�n#��'P��I�ɌVJ�^<�,�׉���֤�?��m���SP��dK��AJ���1�H�P��Q6�	�Ŀ+����+ju�8�����[��7s�/��#�r� �ޑ2q�V��������q�q֩�)G�����K!݂`g�,�\�P$��l��0[ͷ!>��b?�S%�>$#��\���^��x�s��"��=���ZR'Q���ىt�g!������}͊��?���2D���u�n�h���s�w�v�M��Ԫe���!]����y�z��A� ��4�I���~��=��A_��*�=��Vd�\¬��8�.��jIv��mx: ��v�փ(7�E�q�t�,�$����T�pH.���d�K%uZ�E���<���&�(�2�A2O�7��h@8HnnV=Ё�)�k��+W��STݥ��o�@͜�{OP}�2�N*�`o���(Pv��3S��Q�Ə�Ey/|qM���h�ED���`���|��:8ȿ�2t{��s��ӧb�fťm�z��̈́]X��u q����l&NF��(��Q�?��_Pޒj\�I�N��0/���\�د h������o����(:��j5>��9�$�ZI��ma`Wwq1�~~8˽��޾��M�����D�/�p"�A�XG��>at�Ck��O?O����ςj�yw��>�?~�;�[|��g\���a���K�>��#��)(	�C/$)-�Ķ�%��Ð�����̀�H%g&�1��!`����X�⤺}�7�k'�=�*Zv� Mjl>i����Fk�Z,/mO���jJ*w6�{\�bY����)�v�oL�;�j��ه��X��vv^�/>A.��6���(���Y��;�'8�10Z���u�����us�ǜ?�ޞ(e��z2Z�(�~
:����V;V��؃�g�I G��{�P&+��e!� ׅ�"���⯘��9O�D�u�G�K.P����M�:v����#��֚�~��0c����}XF�+�v�9h�6��ow�BЋ24��wz[q���,JlK����=(���K[�����92z1k�?Ņ���bȺQ+z���v��aR��S�����م�-m�	G<�/����%�����WFx��~������p[m�EQ��7H��d�9���"N����n,�ԭ])-5Rb|�����|hk?٦�9H�O�Q�+}�Iz��Q7ǬA;q]]��?��ܫ[<p�ʶ�!����{��r�D�{l/���Rr�jq� 0B7d��Y�\��N�³ŵ�5��s�y":�^<͘�o`g'
��Tv�BáJ9��0�>��g����U�s�H(�$u��&��h# �P7F�V�[��sn��a#K��GN�Jkx��v�Z�	�U)t��7�d���[<�r7��	���Jw����/W]�����eN9���1�����K
��?K�q|e;f�#�0	�;�.A��[8�V�m�:k�gĐ�r,v���?^|��I��/��G6�뜺j&���A���˦X㶡�[��mf�t즹,KVN*W��ʭ�����"�ㄪ�	d	�G�a.���9�R�8U�`�P�1�:zm����R�ۑb��UB�$��h�=�~O��������x�!��+�+d`f�6����X�`���BP�fPq
-'����
�obF*7:x���|�8h�~-Z<-��oi��l�19&��iT-�E��C�X����@^3������vk�E�
��1������PI���{�Ql���R�U�F�Ţ5( h�1 �V��
��ϛ����e3���?�!�؀I�E�k{��]s>�R�~{ f�mmC;��	�_ 2~e��}�(cn��E�hCEE����P��	V�Xc.WRh��V�k�لS?��[��=i<�ҽ�����LU0��"0)���������D�������ƕ�9"��і��&ړ�K�򪫑/��K��1ɷ�k�}�q�i3�N�Qm��4\ɱ��t��n+�w�K�N�XE\��vd*�h'��?�"�k�0�R�d~|����� [<�c00'�����_��*�+�.zM��5d'�����Y �[�"�x��,WF;�Ɛ{ֆ�)����oCP)L�X~����ˌ6ۙH�h�]*��8�qS������?�!����-"4�{hb|/8l.}JH`�{�&rr���#��F�3��[l�1$���D�Y��e���@Ԗ���a���.)�j�>^�X4b|dWd\�������I�i����Lh������,M�p��W�	؁�����S��]���/���45�����ћ�s�V��KWp���!��^��9R`	��;<��BG=?ϸ�vk���Ѿ߬�_J)$�ni��H�pW[I�Lr~[�����T<9?�d5Q��V�A�PCi5@�LZ.���d�w�}�k�ֲn��K�e������P����ԣZR��q\���G���O,��&�BB.s�.���T	����௨ڳ:^���&��R\�Q��KCbD� [=�`oQ��m9ѭ�Է���3Iw���P��7O]� �,�C�Z�8�B �f��S����O��n|��g���ľ����`o�~˪J:e�Ж���{�����CUW�H�HZBB�8�yȟ׍�:Z�6C�YW���.�nO�˻?N�=���rh����15.�멱���l�1�%ۚO�7�T�;���E��bY�b�KgXOA��,�^��y�vJ�QЈY�>���E�9Ƈ�� ��k@����EŶt�G��,E]����n��f\p��B� *Y�D�0�zΣ6u���Õwŉ �L�H�������I�5��Y�è+#��>~����(\�X?��(��(������:��M�����|�JD���&ÂM,#�|F�F�Y��c��>�a��Ps�4�����	P�u%\xS5��e�ա*8���{� _j=R:�p����cQ�M�Z�R`�|y��PfN�D�^%�-:*��c�vr�`m���w�ɓ���ꆅ�)��P�dmca=�5Э���K}~�ڡ�v��DR,����q@���,|�v��+�Km%?t�Ƙ�������C��Qc�@��a�M�A��=	�e�aYss{=R�m?�R�W}��72nh.|{翨�[���C�=�,2:�T�d�r��X�k��A]��m ȿx��$)��=e����z���[�!�o%q�	rq ϟ��\m�*6;�LV����wf���Wb�Tu�%�$v��O5���`F�V���&�^����W�]z�9ߝ㎑�<�-j�3,������ �ʴ�/b���H�{��7b���R`����5����.�-1+`K�u
�j��L>�G�l��=\���(��`P8�ʭ�c���$+�X���[�b�M]�U�y����7�W�!v��>��;����G'�:�������`�]����v~�ݕm��%��ak3�J����,1���3A_3eQ��7�jT�Y��o�[tք ��Չ�!T����U|ڙ{�������^n`��P��7��ZBI�@u[[B�l~��e	�ܟu������#-��A���8Yȥ,�$��3]Țiq.5;�j���(al&?�*/%%*����L<Pu�2`#2UCq'G��_���%ƍ��Ƕ��<WN����8��
�S�GV�����Dgbn��x'�ٙb��r��.A
��������`/,܇W�����WU�Y���i�s)Y�v�+��J�a��T�-e��U���k'����ӻM��* �ء��<_/o��&��ԋ�v&JpN�8Dh���H��	L�F}{=鰘8Y���W��`*#*��&�M/F3��a�
[T��(��E��VH�����p��+>!�}��m�6mv퉢W�� N.���Œ�񍺢�a�x#6���f�ؤ-��� ���ڹ�/{<~~����=߿6[�bl��A����B�`6��zv�f��Kb)X��ك[����\��rM>�M�MY�g���~��<.���
����ŇNӯ��'j�+������8�,�gcO��ܓœ����0G.Q���I~��ܛw�.�fi��*s�;��)���ϼASu�a	/�/w�JY�'>����r��Q��;����>�>��3K�$�Ȅ��le��֭^�H?��j�T�R������ȗP,N3����R��.{Ľ@�ʜ�T�]JlɰQbT_��x%æD�Hw����Jo���@�c�3Tҭ8�����~xaL����{p��.z��N������SP�c��UX�s�\Ҍ��Y�b���ֶ�?(�[$l3�kw���Z�67� !L�I��y�P�ޥ��j�<8�]O qs'�{��� \\��4�����i[[�Td��<���_���W__y��/2��$�A���8TT-�Q��l�ը�ƽ�Ԟe����� �@�}�3�`j�O�^Ȇ[n���-�vs�4�[[K����uv~��^ܝ��7:�3�?Uׂ���G�J��Y~��a��;h�]�->�_	�w����yZ-�ɞ򿶴P-]R'������Г�����M��2Y}_Eb���Y"I��	���Y�ُx咆�B���~��:�b��v�c%JO� ��C��Q_�{���V]I��7��M�ݿµ�5�B��7��3�;��[_�Ca#�V�O�g��ޗ��=}*9�?|�f��
U sV���]�$��\9I��Ҋ����Qӫ���퉵���7x$V(��("W��c��� !E��1[2��7��WP��V�<�8�-�x���5�"��&IDP���ٰ�{��V�,z6�#x�@�م��IyN#��4B�M��J��C��y��҃�j��&�+H.�5\�??֝�hK�o+}���^�s���
`�ٔ�T�MX)�tD�T�4Q]I�5�-�-���%*(�,�R�̱��t�z ��7M����E�����{0 /���i��VVp%��{�~9�⚵l1Õ��#B{��Y�=�SL���ꆆ�6�G����^�}=����`��zae`��5�������Fbaa�A�;�E��
q/N #�T�iu���C%~���9��P��5�gP@RO$��U�j��={�4��U��X�5�3T�:��D?f��t��>��B5h)��L�*�m�$���Y��;�3��[!�V{�����r��o�fB�t&h�7OZ�Ey�JWT'~�������ŋ�)'�"T4=o8�M%ͯu!��.��#XH���4�
Aa���$�֛
�B��+�;�X������"�R�W̟d|U�c��y�آ�e.�|J1����~~��/�"7��}��f�Խ����hex�:�9�q/�(w E̵�,H��5.�p�3'$r����.�P�@��'���I�M�����������B{�#���,mc�>�ZK�/;賈!#�G���uq�Y�1\1�o���w�M��nx8YP?�G�0�����<;1�y����>���e��a�~V��yP�ƃ���&XU|վ� �,��Qq���(#��ah8��2
��������F���\����/5���G<�P~�hTo{>t�Z�K�{���8yt��SnoX���4����;�ɚ�K�l��o��s�Ұ�}�c��Ϥx%gB֋�6ҼS��7��G��L��n�he'��]b���G<���#�o{����UbX������Cb�=���؜<�V��?j.�|s���+���}[��<K��G7���Fa�����d�$C:����}��9����sd��!=�-��G���߃篅Z�X<��d�z=8���?��&�E��X-&#�o�����X���w�L�?"��:z��=��p��(��"64יh�~](=�{��6oPN�+���J��S�`�����Q�q�w��_�~df�"u�_H�?�4)a�f���ۍ=�Z��l7��"��>�����{��v��%L��H W���:�Ύ�����3��6���Ns��fLЮ���=�0�9/�k����~b��W�lw���y���$�}�G�š�D���2�?�{1�pq�y��B��B���U3(k;��(���
F�����3zџ�6%b��A�2VV�2�V�B�&#W�
j��Z� )ޒ29OR�œC~E�9(����2fk˴t�����)����e�L$L�����g�0A�>����Z^�&�,Q�:��;9Mu�#-,��*�_�Pǘ�҈>�[�������,��u��384��U��2������wv���r�5�q+��cɬ�$�?��_��g(���}~��l2;ZQ ILʠ�[��^�8�go�8Q Y�/�GN��</�E�V�w^�ݼz���u"��g%g&G��, �����q���8��y{�������Fp�9��9����4�>][yQ*[Q�_X��<w�4�e��PNH�r�� ��`��
�L0�R�9��vl��A�� J�ܢ`m���x��z�J{��L���aε�m'�#Y΍_�ou�w��mr5�C��ؚ��v����*����"Ɨ�����=�4��u��r\�DT�c�y��UM���h�=+����Nߵ}n������̑ͬ� ��"~dRrX�?�/�S>��ы�>���w|�Q�v�r|�_�^�4�Z��w�ȝm�jm�e3��(}����&o�����҈�`� �W/��6�}f��m���Tn�z�f�P�@�:�qs�������{[�ҥ3�$�|���DC��^�~��+���f�ɼ0V���Y�O-9u_޸��h1@tw���U��?��Zyl����G���_+����#��?c�a�����)��/kH���
���˝?,gΆE��w
R-���%����eY�O��ce&�ZÔ�W�Ҫ>>���:���{?�ʕ�
H�
"ݝ�ݡ�tHw���H��<��K�<t��!�����������u�r��Y�f�g=���}�7��?�U�#����z� H��m�󆬧^�H��QA!(r�1��d��~�8kkMC_��R�k��O*����Tr�#�����i��S���ezm&JG��|!���"��;^��ŵu��ll���]�SO�^��g��((zl�e�w{E6��
��-Sȳ��5taf�p\|�ⷥ
�V���֡���y��Y�J�H���il��,dfCx0��ە	V�pQ�,���&?�j����)~:�8c�s��m�W݀v7���+L�ֿ�6[$J-*��,��p*�zcG���SV��.�T�� ���4F���7n��S26��Ik�]��"�K>v�_P�`�?��i8�%qBz�Xh7�L�sd�FD�?��?��𗏖���\�"\F@�5xy�)�)Z�ԏ�蓸s��:�����l�U�a�Z�gf�]�8�
((pߪ0S��I0�{��f,X�o��s�T��nvo���L�������k���}3:����62�"&���V߁z�`�˦�e�h�Ǐo��0��gze����M+��V���nzci�mw"�j��"T�',ut@�1���R����=��#af+���s���*��dd�ts��.���	�����>���,{`�䉈�`�Q���ά����͒	��(���JlU<�I��p�I��9,�hdl,�-�4��)v�f:�x��_�"k7<xAk�i}��q��飬<􌅏�3�C�(]��&�n:q�Tf�n�͘Do��v��u�[��*j�j}\�%�aw.�?��o�P�ː�`�v���;�Ž����/�7���wT�s���ɧ,Y�,��S��/�z��ra����r �B���vRL��d��[-V�Í� #�Q�ý�ۿ5?��"�q�#�X��x���k+gM��Щwק�y\���_HH\1U'O��n~t��j��B�D��:�N�8��&5���ܪ-����`56c��|�]���&��Z�1��v��m`�$J�y'��lt���}�oZ|�.�	r[/P�y����u�j����ĺ>���@����ɧy&�""ē��!`����<�Ƴ�~��g �ILT���O'���`��"--��`�]1!z�2m ��+�h�����9/��]6��Ĩx�� *�,�kPFF=aH��W�]�Y��B��i��tA��� �Y���W�E{�U��Cd2���iojs_[W�O�D��ah���|����u�gb����v���X߆����q����>������/8��(��Z�� =�����3f��׫PN�����|�1��6Gۥ���N/@T��P�?���G�WK/����
k���)�*-ͷ�F����JK7i糷�����N��8���P)��f	m��J��׏�55_u�(�f�'��6{�)��A��HRS���jb�&��Ng~�`4/�5����[$�T����߭��
����Bڎ-~z�̕ն��w}��BX���Q�%�f�|BMQ�����-T,�]2wND��]|^�#$��#���CLuc���*].�4���D�Ei"]U�x`��*�a� ��iҵ�����y����E	-��ן/M���Mj��X�q���~�*;�$֣�J�����ؔn*��_�����A��mퟭ�(&���3%_�<%=;:�8=ju�_�"�M" �ˮ��)�qYE��:�Mn�By@��z�s��H[�9�U�F�w�O��-�M9ɧ� ��5������J�;/��lg��9׺f�LC�c��ss:@��F3�Y�g@*��1�/w�%��,��n�{8־챎�k�����6�G����Zp������5�N��"�O�u�N9�}uF#��޶i}�m[{U���5�o�\8�+��Ħ�V�4� �i�Y�����Ҧ?ק|�����N΄��ʴK�t���������Q�ƻ����;דEk%%4a�?ț��.i`��4o���}1�1�#��q��.%���cDMM�ԣ>^�ՙ������40��>���C�aN�i���o~钴��A�sS	Co�&#�Z�-A�8J�ač�O�>*(#���j��C��x�7�V'�2�l;�i��>�)�c�|���k�,�ÿg7-����K���T�>IۊOT�JuD"P�#L�u�u��/ �)S=�e�)!ϐ��l0<��k)���P�@��׷n$��G�G;��1sh��<�!o]���7�gbӮ�644���qH��JV4����������=�c��J������cRײ޵\Zz]]Ű;�ށ4�.�^Ѝ�u4Q�oG*⦩ŽCm	((v@�����m?��:���oz��pw	��@��iny�>tl6g8;i��Gs�SPCcF��A��])i<���\�DB[�'S P�^�ah��Vih��eT�qsb{����-j
�J�;=�1�بũ�6��C^0x'���J�))}��^ѫd��K\�Ջd�`e,lLz&�M�i+���ȴ�lߕBx��}���dM���ۀ�v�.�M�仝z�tDa#=^ޏ�.n�/x5�~폧����cVV�����	�ަ���y6s(e������48�CD��=���";���e�j�2��(�x�ὑ���%7�����yǿb'k7�&ܦkq��{3���E�N/F��D��\\��H�dM�1Ǉ�{�ř��wC!@�����r�13�1'���ͣ�g?�#���xz�ķ�Y{��U���q��`�c�,���'<�������!$�ّ܇��z�$��l��ST�'���:��d	�̕��M�X35a���v��H���o!�m/N�S�Ei�&���M���Q�%�ZE��F�|!�f�:��
��p3j|�E��k3�~VP���6iP}~\bS��^����]p�,'ӝ
hY�3zYOϛ=ID��G���To����n������l��GU9s �bVLٟSo��3��.$	���1�ދ�S����8��G�z�Q��bWZ�<G^/@����S$5����=�<c���T�ɠhz�']�(��*��
>^�˯�������sG��ɃS�h���N�Z7M��C��'8_���� �ӕq�'�s�:sҏ��
�孎>�c������st��>�]����>�'6%r��M�%��}2xf�z�0�ut|l ��,�P�%z���7uk�t/:m} ��x�+�(�o}�*���7�]��(]�ס��Ʉ��Y����gM ���bxMVvjw�J4VV
wv����'��4׋�Z��'�ƛĤ?j��\kM���B޵�Mu;򣌌����E~�g�Y�c`w��Ο�&����h	�\�M���#�7�w���`L1
uC#n�4��ŵ/s�&68��g��\��G���ݧ����7T�����>�gp�[f&��긺ҩ�|�}����e%V[QQW��+ۄ0�0�!Ƴ1~�&KC`����x�C��R�P�(������ذ�7�e���'�o���f.:�_�noO���] ~dV�V�^n�3�4Q!�̦���%q��4�E��	Md6/�7�V�tK��W&���N5����m�>��(f12WK/t��a�!�,�:,�G��z�%����Iً��]l�Oӎ�ro<\�C����6 ʟ&x+�D��f��vc�~�:�����!��#�pxWW��/�F윩�H��i�YN�f������[X<�\V`R%[�(��S���x�oi0�L���J �9�/���%�}�ӄ]e2�w�45zo��Ѿ8����6�H��"�s�@A�km�kx̗`��s��&�ussMM�-7nQQ��j����Z)�9�?���R�SnaA�k6Pnx8�������U}kA�P0���ym�
%����ס3Ec�9����F�pm?҄O�߿gX3��K�x�wBln�PC뎶��Z�ZS�h� �;�dV�����5���K!��0ҩ�����Y��eWGHVv28���X�b��\��-$����BM
�C���
��tQ�V=�Sz���L%zF�9{�֠�E�u㮭�>�����޵ڤ=u �DBڡ�C�-+� )����M�@t[S�߄�4E�����U-m�wm�����K�;�1%]�%>�x��㔔b����֭��Iq�/_���m>�ڲF�#r}XQ M��oƃ��{��|�~�4���Q<둷�����]�9"l5cR(�����\Xh�KHPy���AC�['g��^%�eED��'�I��jrT��1���A����ʪs��f;bz:ژ�̱bW�k�}]�Nƙm������*�(9�;� ����/���t�]]�����z��Ø��|�?���*�~��w����j��!Ԓ�q�����΃�i��{�L%�(��	��g��8���S ��,��~�޽cm��ٌ~�3�\�,1�qTMpm�������N�n�v����q��=%^;=��'�n{�*��`�ė��4��U�2�JCm/����-�XJ{Ɓ����Cl�]�'j�OAW2����	�0)��x�ڜg��z��:�Z�֧��Ma0����o��E����������_B2d����%�WE����3�,,�q�ǆ��eJB���03m zr��ԍg����HE@uR���������FCN������7c�Ώ=i)������6�a؇GG�g��6��A�a��1��I�7`Y�@>@w���^��z��Q����0��`���؇}�Y�Vх���@������� t�?q�|6�q��2Z����K��Ig:
D]�%j���0�5ϦWe[ϑqx�1?��?�siܒ���I	{�9� 8Ad�����p�)ҡpr?j���M�,�#ɑ�Tp޻��-��S�:�H��:�d.:��(�Z�)ǧ�Z%���>wˉ*��$� ُ1�#v�q��a���ʢ\�oބ)v`���o�2���6nw,,5#(D�C�l׸n6��-&c��i�''�c`b���$ȏ�~����ɽ�����
g$}�LO�2pX6���o�ު1��b����O�9������=��t�������	aI/{Sm�܍�BC}�֑8H�a��G�LL�X�_Of3e���)�}��;?f?�����8��@�'`,�(w�;�fw`ⲺIڀj���T�������Q�l�����G���좍3��)�]�l0�Ɓ���~�P�����E�7���+��8P�������iZ`c��+���{�D�ғ!a\a��O**Ｖr+�����@��!�n�@�7X	�}������Z��.ۙ�Ok��G,CƧ���ݻ+��.[��e1�a���Z[ZrR�eqAvs��W-0�!"u�<B��m�9���H���ـt�:CR���
;KK��,�66�~{�q�,�Ҙ`�� ��!��7��[�R�h�d�tWܽZ��c�El:��&ꀠN[�\�R �~jh��}Z�`cC�n�	�o0ا��7��[�� ���
&4��6v⺎<s��8У�ʉ�C��~��[	�p��d��ha����X����s^p1 B���d�t�r/_��~�[�^؋�D��'@(U��M��e,�1�9�[a�{t�z�l�RW<�!�/zg'�J@���ߝ��NrnA�jj��<� ��	�/@�z�$R�lu��1��(~;�8�~���!B�h҅@����p���|�&�� ^�{���Q���PѺ��O�;I�_�RP0NcJ���YK���r�hM�&�o��^��NNqPsv�YX���"'�!����k8��jQ�<�]���"ږ��D�����Y���|q��O���r*��m,B.W�n��k�RPsH��u�C"�)�9��V��Y*_�r���&:��m��o����j�F����a�N����ޯ0m��K�l�	��{z	��M����^L�d���Ϝ��M�@��Y�S(@9	��y��zE6r��#-�>4L�5�`��LzZ$�8���Mxr���	���F�n�����/�4�������_�;1����L[��7w�|�=��C1[H�	aJ\�����}C�t�87fFƑ��,�'��j];�s���@7,�i�������0��U��`�f�
������<���ui�1�]pb�����4Q�~ͧ~�]���*�`��8�����	M���&&�޼y���1����ifS��~�����	Mr����b�f0N�N�@H�U���f������j��j���ȕ0,Z-�h����jSJ����aF����eGS����.Jv��>̖�&����$t�����`�� �c�ؾZ_HH(�X���ICCå��BV6�����Q^����5>��ɑdccv�H�����r2)��$����*k�Xpʯ���+���"
5�ճ�˹u'��[����mP���b=I�,��6�}Ի�C�O|68.�?VV�G��1����TU�Q,"��hA�����ma�%5�������Yt'qT�0
���Ԥ|�;66VPT��꺗��WPP O�0�R�b!���zJ��F=�j�a������ ��\Ы18�]]]�b�y���$�ɻ��vuvrQ���t�0��gǱ�Y�n���Q�P:�ZlIf��c��'H����M�/���B�9;�)99�e��,�G��t`���+ꆆi/��]]r�Mp�	iG����)���Uk�4�].�������8�D���ڭ�I6��m�s�������0vKMQ�z2_����.`x36�H G��cK�-$�ov���{qkj%L�D��~�SP���fE҈�<T^9=ڱ
��皆�vn��u�$p7�M��K0��t�и�jmk�D����sWw���X'5�Ez���w��) ���v&zEIŌ�W+;4�!��	�0§�����pP���|.�n�{4��������跎j�zU��K�}+�����l3%2��q���W�&����2Փ�MT 6�g�3S�@�<�ENO��p>��M�ϺJ�+�ؼ��H�$��֖˚�=I�1��e�J/,�k�{���7�݀1�!��P�Ӎ�����Q6��G,ZE?�ͻg�rhD�hOg��f�W�y-���W;dЊY�Z�Id�����|��\���(ˍI�r����k%�<�twȀ�Z�stg�?-yf���~է�r�#�y�k�x-﫪���*�O���[:^]+A��.��+7��:����4N�c��2Z__5�go���̌�pd�b���*��2\�D�en�_���f�
'��Bto}��p�8#߽e�vγL��^�v'�72Xb�%o�lBk`��ۚ��FG:3�3��A���-n����;�~�����M��)�Ì��L�!b�|v�ښ-B�B
e�NM؈aۇ*'ҫ*Җ�4�8���\���;*������쾚r����30F�����1�W�BP���k���������C#�cI��x���S����@>^޼�&#111���ۺ:a��J�0R��'��e�����
J�J~N��yW�h����ᕦXj��l_*�E���w�����U*�us4=&��I�����nյ_�Q@ �B%�s¡A{�,����c+seui�A@`-����	i�r��m)}[^13\��ؾ�B}E���^.*�����j�Q���4	�"S�54]���"NO}��1��a����㴍T���Ђ��[P�ɯ��N��۽�$��k��3��*�o�|��������f���d��pYG����s)0[�ˋ�/,P�H�@zl�L�> ����x}z��}�\��=��E#�M�a,8��\��_T.�����U�Q6�
���#�7��Zw�?����\��*�?pY�������!�b��4|�=�k�� V�{%�||�P������0CA���L@K��),��Cgec��6��dۋ�^��|D`Y��j�7�
�2��H9�x��i�����׭�k�خ�boE��
KIe9V��q�QSV��;���F�v���M����]:��!��b�FG�ͼ���W����i*�����=:z��{���TaLSyCC�жP�2��a�������py���
��t�sO��/.T�'�G�(�B-�ׯ_�Ϸ�������w��v�)���"�Ε�ɂ�y^.��^YYQ�����*����.(���&���;&�{^��2�G��僝E@T��0jI͡�8�Y3�RaU�����$>v�R�8�M�*/?�Ӆ8�M�Ҡ��T�b
��-����㒋c��Ǣ�x���eN��D�_��2N&�4DG�`w%�1�U��
�Yo2	����yC7��p��LA�Tԑ���"��~��
��*BKs�uxd���!Ud6*\�f}���қ�����S�(C�����ӏ>V4;���_F�����y�
y�����AU�N���37�ɚ�~����P�d�j����q��g��K	h�P�y���Y���(���9Ǧ�\�qfxMM� �P��n�N��������т�f΋?��O�i�p�����VT��Ja�
4M/��uO@����ϴoPf��ZH�bA�pI�3��*ױz���{��_�`ym6ޣ���"��H������K4v:��Υ��Hl��d���n����gФ}5��d^��~��C�7�S��G��
�-�7��ͥ����J��jX��rQ_g��T[����M�X,G���8�)|v�=)٧��g�U�w>PPbCBp|<�/��(q{|��V��ׯ��� A
����rPD�T7�!��
�eX���XO�_��G3r����e:
}�'EF��|��ݠ�,�h7�V�L�Ą��jh�X���Ҙ𲏠���Eb������lN���0�Qi���_6�8c~bfa!������⦾�B��˦8����(��� O)`?��>�Y��nd���`�eI��D�s%��l�q�k �OqYJs�ZwK�Ă-�����kj�Hz�̿E�y�f�����3��&ʁΘ{8�C����>�'\b|�+GB�8.!�03�	(�p:̖��oB��'v�
�-�YTP g|q���TG�7�zz �!�镛H `}��܌�?���Oy^���j>wm� g�t-�hM[�Ż��_>�h�M��%d�UN�ؚ���H�0�j�fh����g��h�%�������&(���1f�)�XX� � 7��"�`T��tb?�1!:$��_E��yx�5xX����-o< �"� &Sݛ��v]=v��׍����H};�]澖N{;�l6�j��˰�ݢ��z3(��/�ݻr^�T��\����4������<�8����g�H�U�����#�:o��i��iI]tۜF�xM���L��"�� ,,� �Ud�lt0�N{���,�D����z�++��D��iU�}���qk=er��g�}��rT���e�ڷ��y���#��������gQ@�HO����^�?"��o̅X�j��6ǅ� ���o�w�z�͑�(�b��Pe+͜.
h
��b>�\�Z/ENNXS뎚�����D�U�Va_/(Ύw?�O'�U~Z���ibe�=K�,� a;.E��Ǐ�IHI��jQ���#�e4�?��ԔO 8{˫�xP�L��{	�2�YG�K\�)�6lAJ*���V9��>}z�i�W-��6��g<~����i�������۟[-�d�W�e�V���D�"�21hh������C����C���돍�3��j<~����i`P�� ʀ�0�&z���|��<�BY�ޭ[���.I��X�\�M��-��m �|��ݕ���G��*
J��E���%u%�\l����<f���^:��)��vn!�
l�����vK��Vc4c�rc����c�P�G��tm�fFF?���b��0�����Xh�ޘ)( �F������br�k�'s�4��1b����ΜL���z�~�q;�-���+dU�
(֘1ް?\�C0��I,-e�N��:͞�(G������Qbt��TZSkqDS�z���o�P[Xk��sR�g�[�Jٍ����I̽�_�0Ą>+:h6���:Z�!*����;������""�"q �5����8��:?ZR�~�lim=�|�ݼ�p��yɁsw�"��7Z�-��G����D��U76.ij��o�o(�6K�/��Q��](/���l�����z��{�ߗV5��d������R�N��T�kn.���񕫫��0����Zh�:��Y�X��J�>{�9��2�:^�5-�U����	}	%�>�	y23wi))E�WH�n�)\��濽�;^��ZET+�1�:ν>?ʸ�%?���Ǹ��	�)�8 �ۖ��B �������O�~�@�}`�'�J`����8v��`PL���f����э��`MU�"r���y�k����3���>{��U�,���n��
g!e!�c$��d�,��tg��{:�,1GG!�pH���^EMn��Nax��m�/to�i�������]���{#����7җ�ơL<��y�Q?�����\�`A��V˵5� k��������E.8ն�:����f�`vDѢ@e�;��9��^�x�� �m�Ud��xY���B_�-ÎC����������tS�Tkh�;�(i>Q*m^��nPu�<����[>a�V�����/7>�����'��R���}Fw�$*�C�j���7�K���t���b��{���N�{6����8Y�q�;�+CL��?�Y�TR��|�����f��(�`/�.m�>Tb$��� N��j���ܲ2�M`Õ�N���`@x���v(�M~��o=��wq>s18sq6SXZ�Ӆ
�ұ͘�C�5^bC۱V�����&�5�әа�d��Y2__�㨋CBdeeb$�=`�^���xvÂ��L ��/|]�[�(�<��Y���ٜ������бh�_�&���B��;���hj�i!����ᮮ.Y��~K���Yj�8m�Q����`����	M;i��_�p�Y�a}�y׽am2<�ý�_�y����+���0 \(G*w�p#�-ɳcT3?���{RrIX�,G�tc�뀸���IAA�\�������|6ь֟9�%w���Y	��CF�o]Yِx�b����1���?s��b>倧�o' �T�����L�U�7M�����j�H�-�5Lh���~|Nhhh��OYH�m�H��Tk�����dffJ6��#Y&,z�s\WG�$����s�s��	�`K��I������d`\��T�������[֫wC��]���4�_a4$����s�חnnmi	h�w��hu�H��e>B� )�z.���H�¸yڅ���UA�'4�k\�>r�iiPl�BI��gem��e���'&��6�������5��W�'X��ϟ�N�6��a�X�$�b��?��}�T�Z
22�N�Ceq���B���7_oNi�e9b���ke.�V�~4'�H"�R���6q;dF��=�hA[�0��|��Ȩ�1%���k��U�U��^�4p��z2��l�uμ���pC��gO D����L�0��sa�����~�D�	�@��gJ�4QڍW2-��ӃRӽ��c�8�x�'O�� F�a�;]ԥ��U���~�Ib��ݵS� ����p <k��'nb�[�?\^^^����*�2�\b� �0a_����*�\3e'd��ť�����Q�	"诅Ql��x�{	���{��
B��;��;G�/?;
pP���\4��3�e%%%��t��B]����q3��~t�ۭi?%,v8���{���)!G���*����7�0Um���Z���ƛc�n� ��9&$�c�@�C!���Sx�����^���D�{A��Y"�� S�Y�D�'���a������ ���4�N:r��a/�< M_�_F�sBNcZ�����R���S?���C���s��ǵ."n��̾���U���Kr���B9�t<\2^l���X�F�&$��$<�>�嵵!e�cu}q���"��%�b���v7ɂ�5O�Z4����{)3��.x-nk{�7���'&�ݚ^�Ƅ8�x�U�����.Sw�BG��l�,ڳ���P'/3�� G�$G:]�.�|ц㻓2S�G�í7>����Zб������~�����Y��6MpH?_)9��U I r���812�;U�])J�M9�}�w��ʏ$�����Y3>�ܨ�' eg�����F�m����᡾�Y�_�8�!J�e����z�{3nfS��BCp�,�z�Kޡ�~�}����x�s.�L���m�h��Ú MpPi�D�{�:P$�܁zP ���N�|0��`�0�R@�:厒ϚUw<[��?���Lz��{?x�#_�:/�P�����W�&G���L���#��U�\�X/�Nx?i�4���\�gV��ؙ�� � �b�K,W�cu�+<����P�,��9E��J�d9�c+~�f�	��r�T�_/���%Zx��3NF�����!;\%%������u"!!��͚Va=f��GA�w�f������w��Nh+�=��f�HGGi����7"P��/7��-Dn-���f���V�D��$o�쀁W��P$`������{����N���j�j����|,//w��=���R�'��7�ɽ�5	u5�^n�G�#]W��%�&]�d~����p�v���>�.Ot�.e����?-7T&����*�p�S ��e�%��d*��V�fb"�衆����<`���t0�x5�E/v�m`�}��z�N�+{�[Ǵ�����'��]ó�fpc�T�c�?E++ր I����9�K��2l��w	7&<��+�@�R���p��"�ڇ���޷�g��GDD�M��Z-3o���lZ���&d��R]j�@eNQ�"0��mRr&_=q�X0������M��]n!7��ؐ��,C� ;kn����|{w;(iP�C�Cɦ̎�V��gV�+%����x~||l[����-�
�����Ϯ�C�p�㌋#ګ��4^���h:]��]7�N��k�`�}�g���'(�e"��;�ھ�)�l@j w��h;U�����w�9D�!ݔ}�8���p)�d�s0yв��\��<����ŗ�c��@&������rV�S�I�-���_Ʈ���Y%��=�nhc��p܅;��] ���}�r��� �يv3�1\]C#�d��دyF��ܷ�Hj8��ɑP8eU���KG��%���ۃj�R&��I���@؍���J:����q7{a���b�H_W׀��T���2JspxPY��zU�f-�t~�Bli�����̞ ��� 75�MNIA^�/7�se�&-�=�7G�@�̻]W^��F�OJ1�QC �I��
���6�Ԙ؞���M�������-$Y���R�4Ot�Z���SWV�*�shؒ��f�������1DJL��M���P=-����u�l<�Zw��6�U�����a^n6GV�	yV	2�t�àFeu�S�$�z(�=;�	ZE�"����|���fv �$�%4�T��S�U7�	U�w��A\�@+���~Л�HW#E6��"4�^�#��)���Tfb������c�q)��^� Fj4���99?����\�+���{6�ܳ�bJTo_�0�m�G��UW>L��+i:.��Y���8AO�F��z(n:����D�Bۜh2�,m#϶Q���������u��eR�t����F�p&ӀMFXXXWq�sf��V�P��lEv�����O�ӈC�A�d������F�g��rf=<Mc�"���4bk��*y?:�dխ~���H<�c�f?��g��r�Ƹ�l6 %�ߍ�����NX�}���Zق�Ħ�rh��>������]�\�`�� 
����bd�ç�'쪙P��ݾ�D���lL]���yI�n�KKS��q�хB��{8��a��I��v�:Cc���U���eXnr�� q�u=;W5��?z
}��!Y���w�!�(i�)ׄI{�.TU!��3TYYO�Ϫ�dV�6��aD���ǖ$%$��;4�-��Sm�OO?&�J�с/o�]�O�bK�_�K�o���`�%��D�v��}��io��U��J��GwAS���B1�/�%��k�PHe��Ԅ�)�1
L{Zam��E_:5��0�@ ��E@���M�8/@�W�69�MWid�SX( ��p���w�'#�[2bG4��,K��t~4�����kc1|�F%���U��h^�@ڠ�������u&���\^
.N{��dὊ����7�\�̎�=�g�"�u�Y-�W�l�d/�!�|���w[�C'�>^����%����W��
Ԙ�@,l�J��ز�>��>�]Q� 7)}��puw_]�����΃߀N���k�ȱ�0�U��\�����T���d� �f/i��+g�v�SxT�2V����0?B\�:�:�ڂ-@�KL�����&���i@��7&��4����-9SLh����1�A�?�NZ�*�\��h1�܄����<CӦ[@���́R� Ƕѥ%$���p���Wc���0Q?�m�(<T�*}��ڇx#��%��X��ж����o�"Ĥ�5����Nwy�v�����`ƹK׈<6@z�ڼ��57���h�H�X��3ǆF��-[TG�jI���j��'�&�`:S.Û�A�z]ڏ���d�p@�4l�o0,�\�I�t�/�l��edd��\)B!�z����Pg[�&DB,l���!\Z��;����]�;*D}���D�� �_PP�&���/��}�W;R�rCJHH�I�#M�F�X^>�)��ۯԑ�]�bҷ*X���Z���!uK�0IaD�n����8�I��Z�͝���WD�_u��i��<	
9��j�Zu Î Qq٘��"�¾Ǖ�''��#`��<�U¿�x�Tj��@�lk-��UI+����3��a�h{ۉM��Yw�Ÿox��2!t���jP�2���ܵ��W�/���,z�:eOx,zc�u��g�N��q))������ ���o;�&�^.]������gaIS��WO"�S�,
`W@��'��$��JGR�#�����w���"V���k�&HyC�E )SΊ hVa��l4Yb�
c6 D��f�M�n��/A"���X��C����V:-�ijiQt��CqV?m�g�`^��dQ�l`"y1#�Ճ�}�Hj�
�H�Z�ͨ!qgK��\:ʹ�!����g�� ���������f㓃M��$�Y�z�#|g�/%������׭0���t���� F6M�Y
Z�`)i���Y�B��
�ܪ���yu�ʟ�� �h2� 6q]N�lGe������y�GR��h`<�v��4����IQ��J额����L5��2$��S*)�5,C3=U� ��PS�� y��Op+�خ�H4c�Փ*�������oُ�,��ո�~�hB�i�m�-R(������h�8�urr2d?tw!"���\-�|˪�� �w0p�Ż�%� �2��Tr��LG�&0����M	�� �+,��#9�%�-��lj?~%���ki"��U�5΄�;����n^�u�e� i;y����^�S�%�i�����~>`6�C���Dꖇ����Gǟ���&����3E�����1��� �*>�i��� G^�.����|�2�2'S0J�+C�?/�/�Y�pV�n���v�_�K�q�sV�y�J������N 9^[���.�`��n�D<��x��$�'��22w�!8_u'�p�̥���ӫ�f�
�dA ��_]F�॥*��].�`< ~��=v��MY��tzY�f����r)�H���]�f�Ρv���.nnɑ&�1թe��@<��Ģ?��*]�^�~P,"-��M�Q�DH��X���J��W<��_���!%9@�Tw�K%2�Vڎ2A������TTf,�gc�,<��f[9�VYz]%�իR;;;U��oܸͼ�O,H[��f9g��\\6hZP <:�U7Ӽ;����(䭞�>t� �c�q�����;;��#v��Np�q^T`ӯR Y��ZU��;M�U�@ ��*�݅ˇNrQ�-v����p:�^�����s���A�wǳ���&�����:』��@����ºbAu����r�Ҏ��� �*�$8(����UU+{(cP�p�ħs��Wq�
t���#��:��`�>�f�oH]9?'�\͘t ږ�}p>�٧j�����&�ʡz�󳓽���4Q��6��5�oU@����T�	D�\�4���0�uR�a&�	��ɸH���/NP��o�Z���S�ц6��؀��LB�{D~���am㴷��"u�ʞ_�ep�+0�QE`�ÆQ�����X�=�O> ��o\������D�y1�7U��<`��^���R���61���$�rAhf��� �J�\���e�O 4{�<{{{��Ĺo����T�c�w*����T��g0���_Y���ڝt���,s�3.e$��<�fK�a��fQPRJ7.���l*��|�`zZpy�<9�^[� �Ȕ=U;!�����A��ws�T�W���S��5���P��a���U�8I�^I�/��h��z����H�'��{Y���)A'�GFV:f�������� h?}zF�1J���(�O3.�d-\B�xO��4i{�{D��K%�g�E�н�-6�|� ���c�mcc�x�i0(�
ҁ��b.�q(�:�>���%HV���[�ӧʦ��.0V���܈8���]b-F�s� ĉ��0���A_a��'n)i�H�;�'?��u��5��=+0��T����
�}���5X�߻�HKI#;�V���~"?�<����[��RrE~!4ံ�� 5����\7/���(.-���:ut�{�LS	�B�B��^���Z��m���e�OpZ� IT��@�������+pW�]�c�k��.�保0f@7t���#�+�0�o �����]:�&�C
�	m���z��m. n����X-'��K����?�`%Ҁ=30 �iiR^������'@��r���}e:�*=��Q4�U�@� �J*+��\%�~s���	�����P�k�˖�M����kaD_�E͵�`0��3? ���z�����Rv��m��&�>�|��c��N)�_<�ٸ�&.�jР� _r�R���y���x���J<df��wo���Ս�\�;_E�'���G�YX"����%F��D�����!�t�G�k"�"���I�&
\/5���O��Qk	��d���+({B�X�5q�r�󩤜� ��I�tTkR:��������C���uD�a��*`��4�ϣ���ι��th,a���D0ֺ���q�fh�]�,�]u9�АWR=ĸ�Nx5S�++֗����d��	��KM�W��R�F_���qY�y��0��;;IʙU\)R8�Zae���-@ ��eB�y^~�߂l���2��i$U�Dw/P���������=��pr�Ƀ{�� �=��V�Q����%,<�{E���~��7�J������Pg�Z�%v��H����\JF�|6�P��0E!��q��tŎ[.��$	��N�4.CC.��֠Qn���y��}|���O�~�����9��y������{�ynUK�W\�e~�qgд<Q(�Jm�>�u�*l�m_�7�ZP��������T�K�2׭[BEE�N$h_�Kρ#I�R߁>>Ћ��B=��4��le���*hʷ<���џ;ݯn:���9vz�~j	B����'�����$a-`5>���a�-zkr7@;L��x0��jdA�dB~=u}��Q!����yh���9ՄkW���ĉ�0o�>�ȤCO���t�;�"���&����y>����*�Je;1������U���ח�����9nLK;;;�j�x�t̛�;�74�G������Z>&�3�p\�(�o6�,#뤁�m�腫X\���-���C��;w�wx�"�9]�)E�c�ڶL<�����չ��:c����x{vl����z%��ٞJ��\��Gw���o��p<rd�p�/��q�֎�k���-��-k�a��䗪��]�k�4���ŗ��)��?���U�����\����6J�営O�]_��n��}h����8����Wl|e;G��䦔��̭�5�j<}��V			Vj$���+�G�/�a|x�����<<�kM5��F���Ώ�o
T�k��4�;,(a��T�I�ݠ\�yr�N.-�$$^���|�I�����i�A�,���Q��͏��I�^`�2Ō��̙b�Q���je��:/ΰh�||){@�Jֆ+Q�l����m��*?H�4m��~&a�������!<잙�֘nP5��՜i����;�-@�S
�uOT�����~����G�킮݀H
����v׫�D�hG	��NPK]����Ǐ@i�����k��j\i�3��/ި�>Q��?��[1�jʀ�N-��k͂@<������I�c�~��gi��[����B�Q��{��l��e|���̀�6ī)�I~0�)]�6+|4#�����dw��>15�/D��/f����`�N�_`2R
���X���n�pc����)��g��%�gP[�Q6��!G]�����L	��;�A��б~���L�"�2λ���=�XԠE��|?�������Y��*hlb���o����	����ͧ<,,,����q�/�ӻE���3�q`�ޱ{Z3��)�B�u_�Y6��Hn�)�ۻ� �4��b�!��a�tĂ���p��?�M�w�ML;��W�k~,Y���@h'���e�;�ֳj-M��h��ȝ�u���=�=<8�?�m}`QmԘ��*t�u/f�:Z뺅��I���nwW�{���||]���\ρj�떛�c���
	G��1o� �n��{}~:B��P|��8�ު��E�L7�wz����ܴ���(�|w����Z�Ƌ$)f�ݘ���|0c��FS�{�DO��~#�����N�4ַ���F�\��X�������{��rb!
��S�"�<H]]��W!��\���eL ���:+�{[�=#�%`�c`��|TaT.}�g��u�m��x���OX�Ǘ=++�6�ۛ����c	��D���ߤr�x��ݖ�;�Z��Vx��nMԱ�q}>�
�/��ř/���y)3)��vA���֧'�??�S��v����fw��Y��g�d��wU��w`bT5FݭMA$�a��0�4R2��6A|��;U����	����iԘ�0�,X#��rm�n)zi���3w�+�5W�����68�&V��� 'G���8�S�/�2y�P²v]k+�Ko�vHJ�MZ��+K�i:x%�+Y����l��P�{�\%ti�#g��a3�A��?n����Tp���y�C�i��=�
�ۼ�Y��zfo �oP�3V����M�$t��衉������:Pc���ބ���� k ?/�4<8���S%a?�lVg�Vk���׫"N3���̀�X����l�0,�v�8kS�G�і�1���
�fm��d����w���i��!F�����>�.A!�u�j<�(�li�z�T��o����f���Bb*2��_C��<H�fhĩ�M<:*5P5���%�x|tXWr�8
洯*&E(
���Ғ�7�%�qk��n�&= ��\=W��;��!I�h"ZJ���XF��1ތk������f�"��u��V�� $�-����R���./�m�%�4���l���4Ӧ͖���l���#`P[p�t������?��t�����7#X���K;ԓ�G���}nA���&֙1����g?X��EHa����.�ֻq�_�x�q�Z�G0��I��Ɂ��L��_��>O���	?d;�Mt�5�z����Ih�o��6.)-5J�k��!:<`HZL'(��I?��K|�����̟_���r��:���z�������|���׷�r 6HjDF���zU����]��v�'�P�t�a�/Ͽ�`W�j@�#��n�U>gmzC�/d�>������p�aZ�#����,�3�T�Y����m㭪�=�+#M��F{�_���<���'�2G� I]|�Wi�/�����23��N0N7�9�dR���ۤ�5�րrODIBذ�z��H�pgT���4��Pݲ�w�=9& ڛ�c،9g��"\�[{��	�F�R��mKg���N��ř �$'��C��ήx$��=9�b���~����Fi/����x~y��w5p/��O�=��/�����Ǟep!�[�|O��F��.�� ɭ��J���&-�-�GHu#�BwE�+�x���Rvɱx�t�:�ԓ�N�>��[��79�'���K�� ���i��=��%�nG���~e�m�#�l�ޢv)�������<�V��?��=�3L��T����s��%����X��_�_h��m����U������H�e�֍@�p���ޤ���a]��\�Y۶�"��} ��띷�ɬ�����Ma����)#�	�ؒ	�������S�(���Ɂ�?��=����hT@�ޯo
^�����1ytu�O뉅�z:�@�@�xz��]v�����F�͇,�h����l�����)���o�D-��f3Ŷ��k*�n']�~���ž�r��O�������z��f�d���+�&�C333C�m����j�^�^|�2֚N3�,����0Y$Lk��%A@���[��i�|A!$;p?m�y?5C�# U8��B4p*!;׾����d��6nV�rZs�k��D��N�z��"�g¢�㭿�m��)�H��p^�nˎ@��E���?[%�B����zQ�3[;�1d��|,0)��xUq���SbEK�o�i��A�e��C�M���kG����`�x@Y6�������e��� ��o�8L,�*��8^�{$5#C^D{�qqq�P�D�=r:'<�.k�b',���dp%A@��=�oi���MvQ����qf$j�����~JSt��+^���ic�v���Nң��T #�ۗ�����|�q��x@��P%jߕ��Z/�XQ�?8%��cU��/� ����4&�qG~{��3�و%#�.�09�������p� �T���_ߑ�PIߏ�7 ��,�|NA85��&%o�հ��s��aM��ty�a�`�	-�&�`9�֕X�^�^6�-f"Ȧ�� D��k �<E����[��\�觻JH�ѽ��g�# m
�Ð_�æ%���T-�� qT�N�����qPm�F���)�h�@+�SjBG��L�D":�����4h�'��j$A֞K'
�����:�b \�;M�kDt��)���y�&D{\�dp��82��Bs�vT�Y�"2d��~��Ѧ&vO���`8)��F��Q�+�����vSu� �����8%�L����6�~�~'��[��y�־�0Lu��H�.$�P���Vv�f��a���6�{*��JF�9�%%%�Nt�-�E�n[GZd�yw]*�f���Hϭ3]` ���#8<N��p�AM�)%��cg6�	(���5Lm�J�?zO�l�?u��JZ�����ċ�K3-�z�@5:嗜?�1"���4=I���^G�Z�}�re�8��ͭ>Mg�u��2t�-%�}�ByMښޣ��7�@�=�}pe�&uL7ZU���WA<��v�Sv`�{�Xè��Bw��/4��}d�;�>��hF����"e���p�l�����r�|��0E�	B/e`vvv�Vg�r�B���l�����P����"��草�|Y�fJC-,�Ǳ� ����D�"��c�!��58��6 �<�C7i�|a������/�`b��_w�w���f6:ֺ0$�c�#�9zf{�$���k}H�$�,L/4�p�0�1i.��q�]�t�����dXfbMS�H���K�P���f�5�B6�[y'�e	�����g�,f��gʵ�C �ղzy�j{��� pkTHs��C��Gys�u��x���\��Η�lX��ͧ����!"���i����UE�o�5�>N���Z�S�����Jı%>P���Tv ����t��hJ��p]4��E��ps����C���Tk߹�0E(2�,2��%���W�L�?�%��k�ƖF�U(�#���Pަ�J}�즶���6ѳ�g�usp���ŎR����{����LtEU��Q>���[7G�]>�t���1���Ԫz�n�W�Dӣ�ˣ4��ǁ�1��D�NVh����M*��������;�x�<)RZ�0��U�9=D|O��{���qB�`��v�K�!hP�L�k�ʅƀ�q%�p�%W�I⫯��y6��_��W��œ�s��3��?�֓�1b���Q楼m˴�|�PEt��������r��V���ד��0s�r�n�;���8r�r���F1�C�@*���M�[<�.�����}�~����A~ܢ��^�%ڕ�W	J"�O�:`��D@������s]b*����K��h��=ˊ.N�/���g?��Cc��s���{n��S|���E+�" �"eM1ȕ;�'�U:EC<z��4ʠ�j��G���Y�g=��D�	.P�5ƞ>Fe�YWD���],���ާ�^Y+������e�wYv���=%��J��j͚'���#\Ũg~~a�(�gB%�(���@�Y��:�Ҟ�4 � �}_\���)5��M@5����׷A���:��M�MSPb���c�'3O�T�3B@ CP���-lϲ�̿`�߽{��$:��3���XN�h3@C��D<�+*�n��Â��@
k���ۺ������uw��%�ݗ�*��a!�*��:K|܀��Q�8� ���7�\|#1��?7O��C� <�٤H=�$/��ݻ�vo49X�Xg�9=�l�a�d�a�@���z�8�C��E�6 s�'3-� �[��l�;�1�ז>����"�47��4��a 0��F�>[�r�:��b{�תcT\a�DtY�b��wo|f��b4��˝���C�r;//�A	�O��9�a�\ssX��~:2�+��6D��D���G�Ъ�*@�N���/�0���m�U�{��S vhHw�CE|{�(9,S0Kbo8���2ƶ� ��P�����b���[0�MƑ�RĶ��U�f|��vu2KO�3GJ����6���j��x&m#�4Ӓ��6ޖ	�^�H����)p0�[ f&Y�� r���l�\�EW� ���^��g�3�&��$�����߫�7��� �o�J:���QQL@{�|�u�=>�mYv68r�����u�Ne��t_s{�(�D��n�{�)�}H��gȒ�? �ʂ�s���Q]����K]�Ӻ�T�����Pq���w֓��o���IQ�Ae:��ݚ��X�6�Xr�)��W��N� ������^�gZL+wzoO�*��r�<������z�:�t�D̀��F�.���>s�^�:F�ƫ�X����xl�a���qޢ^�X��X������w�{��Q�ּ�l�LӳȲ���5't��.Dyx+Կ���B�\W���8ݨ�PY��^B�qo�ċ�Iuz(Q�l�N�E�^4ps��8�R�n��l����p-�f�K�UXd�S= �h��8��,L)8T���6?5:(���n�����!��<�����j�THπ���F��aZ��[�	�<z��퍶 ކf3|<H��E��G�n$�>G�^񡟵�F�`x�F��g����UW��8��ڂ[��S	?�{� c}���ފ���6��耦���.j5�gu��B�q�`�&��CfŖaU�T7�ܪ*��b��]�����M7�$7��v�8���$QU�f�H5y�Rrh��r�ʩ��p���zFi{_	�Q�)^^�Cb�תj�W��! ��#k�X���v�d@iL~��4�P\h
�&�Y��)M?M"�iw.'�0�DD���,�l���ۤ��Ε�P�8����o�nP�¾X|J��Z��R�6�hf��_6p?��I��Vn���qV)�.�w�ɽ�Z%��(_k&�<l!�����JJ<l�[��Q?�[����^%l#4�yckʞ�X ��	NjYHX缤F��p]���	�����9�TA+�� �	u��l��f���}X���(��\�N����ﱹ1\`��m�B7ܰ��6��BGu��YL��YG��$��d�9�D���"ZQ�kN�/���^�ޭ}nmC�#�~�#�T�.fж4"�]$O�y�����H",s�]�F���F�Z;�(�f��[�2�qkM�����g�P�L��_�Y+nhF&���PP��\2��+�ˣ���R����ˋ������$[�z�O<wtM�H�GͲ��$��� �A�r�ڳ�X��@�X2��C�^�nBT�+T&�/V��^�H����1�4?�6KӉ���z����16Pm�F���Ȭ��^�,*$��F���C�գgiX�u]>�~"@#���>k�XM���k��l�B�}�=��2�[�h�d`��3T��C��y,9���
Iq
��B�n���XyU!�=��Ç�i����H�<�#�n�:"��MM���s8�"_��O:ף�L��1�)�����K�{�f_�OF#c��/
r�����7�to"�j�������m��Qdi�E�1��J���Z]m��^y�o�$�t���vA�@���; �
�x���1�<(�S�A!��k~w��B;E�y=�J��%6q��Gp׬r�B�2v�Ad��z�#��˗HZ�:`��h�!;ۺ��:�?
,�4x���˙|�Y�<�f8�kU<#���?{@u�A A�����;2�R�1�/5wv�!��~˞��36�@[KK��d�**E��-aD�N$�/S�t� ��gFz+D$�.
0^���4T��p��xf�,(���Pp��J��D8��7�7��}?^@���Y E��+ZZT�y� ʯi�K��h��ݤ,Jz��V��}{���5$ii��D[yh�z@�m�
p�z`(�eߟ�2�z�<�jI%�kjf&M��M��	�X��� ܻݎ8��
��w��L�A�>SI�ƚD7;Ga4ĩ�m5�:C�1��7���{�͝�s�WwW���~�b93�.+z=�b* �=���	D����g������R"~v�_�UAL�b���E�tefnTV�)�Exn�I�sa;��;����'��r����,ڤD���莽����{��B��bM��E������ͷ��<*Hx%P��3B���V"fv"��:�ȩ�ɎT�&��@�kzфR�C,"���JE���(7�<����8:���T�6���k��X�}j��,Rh�,�G���t���H��w��0������2�ت�v�#�>���,z!RFh��������/z�}�e�@/�����>�^�+1�6�.0��xt��aY%a�%CS�ʾ�5��~�B��������Q=-�T0��>������D�oP<��m?Z
�Fx�����R�i?��Aɋq���PJb�Ж�c��],�Щ�R����l�*�^ҟ��s��2����u1�PE�.Mӵo���3�r�LFcSK�sI��b��Eӱ���חP��טR����0��X���JIN�����w���h�O�;ԋ�<��w��e�s���_�%i�ϊhg�����Oi��%��Ֆ]�]��$����=������LM52�H����y�?�6j(��;��4�	lVV�"��+c�;-��P�b����x�L��D��V�]�8��`�!����̿���Wↂc��Ҹ��Ǐέ�,L3|v������Dt�ɔ M��a�S۵��������v|�]�ˏ�ʊ�����h�J2�j�akב��&�G����U��������g�y���ܿ&�e�]���L��b��N��h�ΤY` ��!���	�Zh!���b-�#��ha��2�k��\�~�3+�*�ٿ��Y��SC���)ş��in";4�J��B���t|(�9#)g�Ŕ�!���˳aۃ�Y��zʗh�c��d�(�L����L#n�ସ��� �Ss��/dE-\ʊł�CS<o��{ Mw��Fve�o����9K	p,W����EQ0�dE����Y5��]� ���+������J��k2:�$N����xֽ�_�ѡ��ʓ����E�su�_�r'��ؤՖ�� NM���R���
�Z�O߹�H	��`�$���Xmz͕�A	�"$�9Z��	V�� ���MJ��<����JT�y��gJ�ɝ}4����^�%�eZ�`ْu먹�D������-���G'ĺ�jyê�V{Ck�l�Ձn�����E���!��w+��<xu����(��,9	��{i��ּJ�<�͔j���\5Z�d���7Z��N������X��<�~�r��o��"�0�q�bb݂a����
����˂�*E"
�M��&:w[�R�e���>ǥi{q�T-�=�I�����(��[{�wq�%~B�+Re��Y�g��� �zF����I~��H�i�7u,;�",Z,p!Mse��P̩&�&4��.*���<c_]�HR4`+I0�	�gkx~��vء!O75�W!�W�滫���"��G���:���9���
�ת��W��>@YO�(";��+����^���w}�ʃ7��a�i�W�Ȥ%U�8J����e�$�=T��V���;y�jy�&̻����K�Oٌ���<����P���u����l]�W���L�L:���r�m�Ef%��#)�$.��=$n�{�:����V�������vp�4M�C]�3∙2rY�Rin��C�ݸ���w�0-q���=�Oۮ8P82}���E�i���O�M�Iޫ�,Z���W��	��J�	��u�T�,gSj�x��CK���'7�/�5��\����sw��h�O%�$���MO�i59p��i}/n�i�3�4Y+�"2��P��x��L�+0c������p[WX�,�W��㭶c��F���L����5�r��dVN�f߽(s��E��M�
��b�SVFj��Wz
����6��9c&\р�SN��ۡKK�t�.N#��_�o����(�i��W؞��>��2�!���L7wa$�f	ۻ�6q'�Ӓ�^�S����k�]¶j-�4�=��@��ǲ��x
��Gg��5��,+���%_y�FT:�n�����7��\���1��)%�t[�rlW�ݞt���X��3�\h;��q~�[|Oא1��ZC��0�s}Տ	�>GO,{B��-�b����5��������n�W֜�������.�e�#���PK   x~�Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   w~�X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   x~�X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   w~�X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   x~�X0%�a�  �  /   images/d63f6a48-eabb-43c6-9b21-e1ae45e934ae.png�v�PNG

   IHDR   d   p   ���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��]yp�U�?�%��+$��@  �#K@Y��(K9�(xS�P�yj����y��M	5�8��c,�Ae�Dd�dM�da	�		ٻ{��~}�i���kz��Wu+I/�ι���߹F�!6m�D%�����<����𶎇��L�����)PX�bS���l���gy�8��9��c,�j_��S�X�V���G�}����!�V����, ��_�a�ЀM��^G0��.P�@�>�K/�DK�,��:���n9z�(���?�O<A�����l.��>++�������tF i�]�zu�k���-::���A�|]�8I]QQQ��O?M!��/������ͭ3�LULg��^LU��_��ԩS�̇' �e<,�>ԑ@L<��x��Ԋ?�����(o�� 4���[�<?�ǂ��c!�6������<��f�������|R��@ ��<�R�������J P-cu�W��B(/��P�a|��ꂯ1����P�jn����s�"�"al���ۜ3PϞ=)!!��z=���] �*u���B���b� s�"���)Ua�F�:u*=��3���,��B���mnn��W�Ү]�����j��CS�3��Ij������K�ҠA�����,�����]p'�b�@�7o�ݻw�}�����	��@������P�.h�&~������@��易�ڞ�'Ґ!C�
���%�"���OZ����μy�(??��ܹ��s���&L� .�F��y�&UUU������w��[���
�wcc#�&x���|'&&��ג��hԨQ�g���_U ݺu��ݻ�������o������އ�yꩧh�̙"����^���'�v�����i���4k�,1w�������] ��X	�*�����V�Z%����,z���ĉt��m���zA�ٳg��Cu�@w�ޥ5k�PAA��LlYY�x��8t����W^�ޙo����X��
����{���|@%%%���G�G�&��,L��Dmm���o�A"JE`.Z[[�"D�
A̘1�z��A_|��:u��cA~�ᇴ|�r�۷�&�5%X��!��{�Ə/ŀ���a�A�d�⫯����6�x��`��;\&|���b��v7��Zp���Ǝ+�1&f>Gm���?�@�9�����߀��;w��eĨN�w��N+���gEE}��'b����'"*���H��p��yaSC໨�H�	+0O�DKxQ�;�;wN�^��~�# m8t���(q?�!T��!�#���,���O9994b��r���#�q�v�g��
 ���Hg��`�0:���ќ{EC 5���B�C1�\���;�%�&�O�>_�*�v��"��b���"��	�h��ի��X8w-@�9lذ��C�7�8�Θ(G���ȑ#5	���T�͙3�V�X�������"�o�fӉ����&P����-`�Ϟ=[��Z���ӧa���ՠ٩#�Z�p!�[׹�T��5mڴ��?�V=eƍF������DY����nb��?�X#�=mz��������M�-��?��S�q̘1"y�j4����N�<Y8+�P�t�S�X%`��`���d��ޥ��*JK��ؿ��`#D����(|�
I55qTV�̡g
'w1B���#�v�2�\��>{�L$3�!h�� �k"�����Ι3g��ŋ���H�����T�Y�k67�C��~���w�f�)M��\=���6�ň�j��T�F_a�X(I��zq��NMM���o$���Sd�|�LA3<�(=�9␙�&̒�x���π�1��y"�ғO^�Yo�
L&�j:�k2��{������N��eb���P~~6]�ԗ!̟V���pCc$�me$��<wT�{��
Xr�q!O#)��_�"=�kZ=*L2rJ��r����Ѓ�V��9m�������;���81��^��k�1�Pg�!oT"��}�q�p����F7�{a�H� �H��y�뵤<��0��M�V�{P)���_��bz 8=����#loґ##��1�~p���Fi�7 ս{M�r�����I��2�n����?:���}hQ)��l&)V �LI���{s��$k6a�F@��n����R��]n���IĪ.���%x��i�O�} ���G4z��qzq���:���O��g.�������J�f��u�C���	��!`����[< n!)��	��� ��>�;ڽ{�](�є�>#5�Bh�"鼫x\��}9)8�ԃH	H��v��櫛G>�3*A4u��N=�Y6&^
;8��Y�����C��@۶mS���_��2Y6�0�'Ru��K��0$��k�ES@hܽ{�ߩ�@�7��z��N8?��@�'��i�#�@h0�*��?	
A9$:���e��{�
�9@hA2����=D�ś�cw�@P$4���G=Ў"w(x Z��fL+h�ǎ���\C�(Y�\� [�`J(� ����<���9����%~����R2��A&^JJY$� �@r��9;��Ξ}�k	c�5�hl�ר�L�DJ-*XڲH����R�x1��ѡ��Aޑ�RM�ɰ�z�@���!�@#J,6����PUU�W�jңG9��v���+)���t�5;�L&���g�r��H	}��tVq��A�sUO�������(=[Eu���k�T ���	!!UV)#���Fr�u�B5kF���*ԏmLC ���f�u)����,���������ه�ॾ�H����s���㸧�+��B&S3g�M,�h�CDD3�����b{�F�`(�t��*)i�#b���v$7��
>���1���B��6*+�#�ʊ~����0�6XK����@r��K@"�s*�(;C�UJk�����>+��Gy�=�өAx�=�6�^D&��W[�̝B���+���bϰ7
��g��b46F���Jc���B	q!��6#57���ۊ��5���bW�� ��	Mqz�%(q㆑�DlE%��33/�^�A�!��2�]�		w3w���11
j45�91Q�nAwuu���W;Q$|�^���R�=�`0Sqq��Hq���`�A���7��[Ϭ4���2�nu��
��F��t��9�r����o<3�M���X V����A&��m���h��h���l��3I�{WOgΘ�l�Q߾����أ����-,�b�TPb�I<z�`$=�|p�b!�)#��#���<xk�C�o��1���9����D�GGӶmQ4qb#����@;��S
�C�D�ي��W3��_�h�2/^�KcǞe�DӖ-�}{,�����hǎX�<�e���c�lA�7w�ۂa��ł��4`@��7Є	��kW+��fv��8w.���ihGll�����nPZ�$���!��i����h��xz�*�����u�O�!�1#�N�"*�|4��e>0v�Z&]�T&���K�����>�(�^{���K`�IC�^Ѐ��j�Д)x�z0]���a؂i�;b��G����~�3+�?��yI#���I��_WSL��R_��>H�&�ڌ#���t��0��Z�w��t�j�gO.͝��~��n��;�ٿ��ʕ)�dI��៮s�n�h��D*)1�&��T���r�;�0�EV��z>D	�kk�٩��9s�c!��{�ݢ�b#��n2͟_ǫ��|�c�"i��8NPd2��ޫ��>t��*/���߰�3�`-/�n��	�Z����xݹ��5kٌE���Nû���m��O��ڊr�1uj6���f�I
蓸�w�++�iӦI՜�e�tlB Gc���A����@ޣ�=ό�<����+R8q�'��JV7n����3�>���`~N�v[�N�I�����?�q�
[D	|Ϟh�#)'��F�h�-��l6���uTU��M8}���������#8ߘȟ���/��^�l1�I�D7���?�z��A��I,�}�j	MN����E��-2�*ҽ;6����&�=p�>���l�B ����c鴭�v����ӏ23�rn�)��I��S�}�!h�"���},.��,胢�����B��ݩ�l��7�-:K�O�ŋw	O�F=_KG7o���u���	 w$�B6��V����{Qzz.��9��m�����&�!�t���"O@Ϩ#G��^�h+�������vEZ���ٰXt�?���^�ԧ��^���
�N��t�	�+T�ɑYe(+f*���ù�P���#a�Ţ-`�5� ����'��ˆ�h8n�8��R��	 ��e����`JKKEo�g�}�^|�E�M��_C�t9*.N�I�AQQ�h��J�7�7yT�9k+���bgB��5�fēٜʂȤ�螬����/X����IF�{�>�>(@c��6�h��]	ū��}�v���/��0�=+c�Ν5��EўGY��$|O��JG�Ѐ�.��5L04�ZX�Z���:z=�u����Si��v�o�ʶS�W��������hu�V�h&�~�z�t�qe��&��ӧOa����/���8]��tխ�رCh���]T�CY�PL4lT�mx��
�V����ضm���rqtL3���Q"�333EWR-|kj5� ��� 
B@#/�v: 5F�5�b<���O_6̆f㌐o��F�y�����@�L�+@(8���:xECd3�7nA��a�#��V��3�ތhj���7h_�a�`�� _z��5q���;[�� @(��������OQ�0�����q_XX(&'C��4��p�
|���T�&G%��
��a���"�NG@xh	��@3h���8�	#--��qGjp�������u$�j}l����|KGP�35hj5��u<����N ͠]k�w	|�Y#�֌��\�PDw:t(��Q����ך�����
GxE ��H$D�е g�i=�,X �A;x@���+̙��Қ��>"���8!g	ųC$d�u��u�R�3@��!�quD�l%�d�Z�v����g�`I��B�`I��l�2q�$�w@v�x����_G�3ՠ*Ԡ���/Gۏ��ԧN�<)N���"�G����;i�$�Ն�0$�4�D��^�%'9J%(��T6�~��K�� U��q#3G�g�ʓ�1�8�U^���vZ���{�xA�N�L�"NF@��H��<�j�� ��<�9�޽Ad[��0/yN8#2��L:6���A6���Cc`��C��������`;í@P4ۼy3-X�@U�9��� ���;h����;�!�7x���܈Bq�#��X�
��<h�q�ƍ�boC +Hi��ڧ<(jV(��*��Pc����&Q���{;��<VJ������PP�)y��K �+��أ���8��F���������;�g������.������/���V�"���_&�m�����#����/�>)N���C�F������M�G/S{��j��<�R�����2�f�%%&��:�/�ӊKJ��աkq��^�rrr&����<K��`��\.,���	�����{>�ߺ�Pg��ڇG@B9e��?p��������Z�a�Ql�	�� %���կ��0u�����͙={��Y���
|J��G;f6D��b���6��(���ŋ)5-����m޼9|�������|J�O�������q���w��ʾU7-GanQ��5��NF�@���G��t��    IEND�B`�PK   x~�X�tԿI� � /   images/d8a77cc3-1409-488f-923b-bd8c8826a526.png\|TU��������)�F�Cii�ii���݇�8�t��w��ｌ�a��g�Ssε�&\EI���ɾS�����/p>�����YRN	��F2~Gv���Qt�\0=�j����.�\>ٛ��9������,�M����,ҡ"$ �k��;	5��#�����,�ڪX^��T���kJ��ޖ�6��2%�4���kk3�2,n�B'x�����H��J G'4�t)6��4D���Ȭ�3~�_.w�Z&���1!!�;�8�F��:UW���,�a�����`�1�m�s�y��>��K�*�oZ�����y���0�����A��U\��0�H�H������a��h��Aa��ڰ1*{�h�������A�
����,��,� �>�4f���,��+*|��o~���d'}T�3A5�*T�p�;d4�qԷ� *P/At��ݣ��YÍ Co4N��{�-z泐�d�J��'�-�҆l�!�/�����|>|���x0N׭��L��Rn�lt.p�r}͛N:O�j����#���AT5�Y��'�7*d��v��宦���ڐ��Uhr����J���e�j'���p~�7<�#�`L��p�a^I AK�꠸���	�����&oQ��F@�ȰK�.��Yɱ�E�����O���K����ֺ���(B���h7��M-�U*������A^�8�E�� �d��I*��t$9܇B�k������m�ڹlt;��=�u��`��C�ל7��1�l��`zz��C'��РQ}�y��ֈ�����_���!<�vۇ�7c.O������~D����|�}~��̝����1�Δ�]����Cp�g�0���7& or��л��w���Uy���,eIA������6��^���zr�_�K���X<x}���ޱ�'�A������y�஢�A�v��U٤z�4�/�l2���� ~`� D s�6т�I��	��l��\���x�t���y�$�� �#�M�����-��$o�ݢ�?���.nEq!-zo���t��؛�G�9�:�
ӧ�0v<G]��=ho�x�����~(/d��j��&�-Y^شG���#�����B迚Fj�(p]�v�'�R�i���lt�aBh3L���=p,�h5�z<������u�����3�W�eԷ���j�*�^��Ӎ���d���6^v��gr�n�{��˸]��'�\���k6��b3��V AG��c��D`�<R�@შY�;4��7�[/[!J�twQ������}n�<p�Ɗ;��s�Z+Z2aN��Db�� &���N�|��d&g��2r?�Yh�[��T�ϣ.�g�hf@�Nv���P<�K'�5�q�����������!��.�*_��%}Ŷ�e���o���
�X�[e�&	'a2yl�iV�4���2��Ql�x�Xm$�Q ��İ�TP�`�[/����[��s���Ȳ�OC[��Z�������������TlDw��a%�miǅ~�s!��./�O�S�k��ū���I`�l�kN��*f�T�J�gk�1�p��;!$�h_�l�2�!�}6f�L�3D������E��@����V@SM7��-�����Q$a�WZ��ͽ�c�I�=S�t?]�L<�	�a!G���I�ε��g�k\���/�w�>ͱ������_�e@f�������o���6�ez�j3�7��4��4zc�~�Y W� Mw�~Hf�������wj3��3*v���?`!W�8�B�f��6W��������=����w8˳��[�"_�_��>�j��Y���V!5�TIP^^�G������R5K�,BL/���P����Q��W9��� N�����O�@�{�f�^	0C�v��A� YC�k�������o�C�Ht?n������R�L/5�(L[�K�
%h���a��9��Kb��@!��[����*�ʧ%sH�J�����Q��s�D�̦|	B�{���@y�/��`U�R�f�(@|L��
��)7*�]���T�a��G��(��p���3\##�Uo�Ux�@��y�!�TKNf9ĉ �����{�r ��}�o�0�xy݊��R2dvc�о�Bo�Ɨ�?܏q�Ji�w�g(��8 ��R����"�ߎ|;P�Hɡ.Y�~m�QuS�	Y�N�Np|��J�Y�_'긋ޞB�	��T��*$�_�	����졚�T�?�f�z�{�r*��ȴ�;#��˴6���f���䢱j���W>�͍�'��XC�H��c�fo�I��%�݄-ѳ��5t��hv��b�M���[�u\��Ii��ttI��t�ѻ��<�R�@��P�ͤ���Z���*�e�����*?Յ��hż���W=���L���$ӶN�)��w����U��(�g��>��7P�^]A�κYs��l�}�qV�a���z����q�����/���V�a����ʵ�7|\җ��d����Mϒޣ9E� {�CLe����tmh׾�d���u{�A��Z��W=����c��%C����@���p��W;ExБ�Y�.ʎgr:ղ���R�H8����#]�-�*�����3.(!�#9����߭O�8N�0#��4����q�g_6�	�fYz��WH���t~�+�?�2��́c �LX�Hc��Ῑ�����\��怺�/;�/��%��Ѝ��~�Ԇ�w,cb&;G��	���ǰ�X�/���@)���ޞ�'EV��N��*;���QζsO��h[��Ǒ��<$�7���Y�6��]�1����/�l������jڜs�T{k���~��5<;��v_:���m����+��I#���d��ڝ��l��WYÆ���a!���؅��j�|y�����V��Vy�z�	ْ1����nm��_LS��G3]۝1<Y�v	w�yuO�,��˧X9c����o
�M�BV[>��c���[��ʙ%����t~����.��VV�'�2I`q[��z��;���y�uY����M
Z3d�j�D��;ӻ�����Y��Gr.}�"�'VCf`�%��(V��̙�\��,�u3|�P`^��ʢ���V��L�2~����^ޗ��HuЪL%�M�O�ܜ��5L��t����q�V�(�pd)��W4�y8�Z$5�#RE����p��z8�\q�{���A+_��e����p��bEH���NA
��	!��Ю�j�Nw�a]B�o_�f��yd*�
;�T 8��虷�7��PگBH�5ٷ���V�	�`bC+�m�DŜ<�2�%PiX?E�j=�&�������tK��V�:l�ͫ笷�p�� �S��_O��o���A@��S=g�:6C�9M��#4�"�u���&�����UW���Z�Lb��p0���֫����~y5bg��D��`t=���O��7*��̚ �7��~��+�U�xm���>���������K�F���>G7�!�0���h�:s���3���Z<�"�u,j������-���Z�bD�2���)c<}ٯ�yĮܒ����P>Z����qY�$�g�*�;��QC��r�rQ�Wl��|}���*
aި<����s�)���Z!�A��o�ӞxI�U~IH�� |�;�.o�	D�������M�"�����������������������Z����R��񭲏JWJ/�/;��Zl�'�����5c'��=���WYlo�U�8ס?�G�(ZE!G&���=�<G��M��z�ǀq�"�>t���6�ڻ*dZ��.ܙ&����O~@Gs퍨�6�$�?>!�;�����+�Ҽ����1A̹��[n�q���r�K�#rs��D-r���3~��`&E���J>bJn3�Eh�o���#�hާ �ú�f��!��HٽD�s9��E~�,�duA2��sp�!���ip�\+F�Q,��mLgz����e{a������C��XQ9�&h���ee9�y]�_(d�NbN���"{T�-��>�M22�u�^+S��
��ګ��NG_&7-��J�%2��S�6������e,`����������b!���ё�,B���ƚia�!�����4�����W�r�-��Fz��}e5��NtH��L�Ȅ������3ȝ��p:	�b����i\
�_��r�v�wd��-��Ц�Õ�}b�7���cYN.n����d�t֪��'��g��e{98�^�9�n;����T����g��q�)���D�v��}3T�A.�3^�gp�U�j�c�����u�f-�ƈ_SjY�#��¯4�'�(֟�_y-R�K�u'�iZ�,��Tp�oC�x��Wub�K��:������j�R���#�Ĵ�&�ܹ��+�" �i�O����j�j��nG�d`�)/�T���+�̮ӆa�i��$��u�zv#>Xz`QP���V}8�A���R�t�#�1�Cw�OA��	�/`b���6G͘G�+T2V�ID�x����=c�uN�|L�:��<2D��X���^歯�v譱�g&����~a|�<�6O٦9�z ?�zm�Q�u�d;�-c\|�?^aXhgK���m>�-��4H��V!'݁=����LȕS��>/��d�����"��6�=[�3�\��M4mgf��n�/��υM 6�J>�G�Zd����g)�pp��^�]|��2�s��v���l���]Yy*��<zCDt��n!�+eWM�8F8q�V��O����C��82�-sB|`��M��C`pm���_E&^|�L�Oyo�No6�;oU�h}&�z�~C7�B��J�Ǚ�Vk��S_�����ԫ�;^��H�1��v��)��hI����k �Cc"�}J��:��m�BG��
$�J��+�$GY�1'����g��?L�ٕ���=���숡Q��QC ���M>;[�B�Z���AB�x��"w���{�!���({�l{z���j�"�h�\5S�tw��@L����T�q��&���o�ժ���"�	��*�(����+)O���ߞNn҂�D?���A,)x�����2%��{�՟�T�3L��%��T���[g9���ϭ�a�������ٟ��z�N\� ���:9;m�����k`��U���E���e��C�ʶ�['���Qg��!��	���Y�aK7���@�#��4�R50����cJu�P���g7�H�C��%�b�^�_z�����=�^#��;��L��bXv�f�?�t���2���g0�Q�K��,�RP/�59I����)�}c��LuF֨ �ܱzb�l6��݌��k�؁���ƺ%� )�ݤ5!_�����h�Q�������<�GWX5LF�l ��
��
W�� -���XZ� M+��[kn%��Ɉ��cy���ɣ��SHJQ<Z�N��h�o��"LF9w��%M��#"��	�&}���Ḣ�����Y���\(h���g�\=��8�8���A .�Y��&k�D&�W5�u�w
�.|�D��׆&Þ�Z(_��Ƞ�t�8A�/S�!>{O��V��g1�������&o�H�\]��6����d+���4?>̩T�(a�&�QD���G,��p��m���Hrq�����k6��7�z�y���w �1rN������m*�S���Ǽ@9�=;�� w�5���	b��<9		m��3�c6�D��#S�GK���q�Qx�������f�� ��J��6��U��HQ�ފ9��ӄK���cK���@7�-���g��D78�k��e���|A�G��� L��E�մ����$�(��c�T{�F��N�"\�����v���1��My�ߨ�*�h�.?�<(-����I��� ��-mN7;<�Ɣ:�d�UO��ʞ��d��ѽ������ZK�B�D��p��~�gs�ñ����϶������c�Iq@�����W���8������W�<^Gf-cɗ��RS1�����/�P��F�H�����eE;݂�4��jh����ۼWaU�L�VtG:���m2��kΙ�|wk3�_UWo��=�������=uɧ�;C��&k\T�k���/���2�������7C�sw���[�l��
�﯇	��$]���I�	r&���rߪ���F¼(��1�͔��Y$���}B��~D�+��8S{��رa�.nn��:��f/�B�Dv=p��#��M��2*6*�0�h ��O�(���9�e�#.�����~��e��id�I��.v;�U�n�ܟV�Ɛ�9�ˊU:p��73T��⋔�	�07�"�Q�Iv]�=������W��a�Y?�o|�fo��㫌ez�D�/ݹ��]�jOiWe����b<���Ҁ��6�'�8r9M][*~m��r�D4�:r�<���"8���ge#���c�T͌n�j_�╮v�˃w9���q�� [��ÖA6o��UR7�n��xiF�Rq�p�hp$w=�4���+��"��7�	�^d��>�9�wC�M���Fzf��V;�}Yf�|����X�R�]Z��	��=�a����q[���kz��1o֍�t�OЭ�W�7º�ER�z�Bn��h���8U� � }���D�7+Jj��+C�%"����@��$i9�.ҹ���h-�`�
�b!WP�2�����4�b%��q�J4\���C9����t§[� ɕ[��LK��l�ì&��eF�k%-��u�&���kl7�|�b��;u��04��%���X��4zU�W�q��8�h�ыJu\b�'u2#�I{3�d��q'�2�X�`l��(>1q��7�+$��|����߷'��`sO����xC5?Ep^�� </?�?N!��jk	X󂬁E4�C%&/q'�}�	�a�p��7�5EOb@�høe�O��/��*0��=.U2)U��N������ �t�Ю��#���ĺR�������b�|%�E,��C���%.w�^���[���2
�	8T`	�V1sR"����ҊzPE�%�:*��y��96S��G�>�w��~�n=_�;�	-h��o��_�M�+����
NiQ$����
�"�l~O�fv�l�M�����)q�I-7�VhL�x���9����mR��U-���4!�mxv����u��谢xǪ)4!����R������(�NĴ��5nh7�ʟ���
�m����|����GO\����H|n�P�g1pLWH��l��]%2��@�U�{ﴪ�j������.�sE�u#JF�\oW����s���0��W/���v��Vh|����z�E����ڵ��~��L���X���y��^
�����fn< ]d5�	��i >����l"[�OʓKwT>�"��[sLk]B��h)Rq^�����~h��8}W�� Qm��dj-����M���\H�}��5��>u-�~x��K�k\��Ǡ		$L:u��S`�p�
wp����_q�#TBϩğ3� ���̵Z5�G�W�$�T��<&�z�h���k�6�f}�������V7���ٓ]R�z�x@<�=.�!qnN�dx8i� ����{X�1@�5�U\JxȚ�"i�;81*&l�h������n�-����N�L7��������ʔ,i�!��E���%��"�h�I�i�z�.;U������+u���>3�(p�e�u��u������ ��wn���j�$���"�d����� �����Z$�� m���@�}�y�0��gzA�>y�/PP�[<w���01[�7.��ooċ�*%�c�|9��T#Pn6PX�lKq=1�m\4�]�tN)%[m �ԉ�Z4�a��O+"6i|_0����N�����b��9�:����vx:,��\O=QJq}���h��;�X�O�l�D��ZĜ��V3�x���s�����K�3�J�	�	�\'~)k��M�$�f���~��l;�dG�㼬m_G��C?�k�,�#,aO~��h�Vˬ~�^���fi�|-7�Jnpv6\��k�,���-���;k��yq�@0�ѽ�/�����#�O_l̒��ܦ����K���G�-�'��	�o
�ft@n4X�|�fؙ_��Zn:�ٟ;<���-.}-�F���v���R��Z��n>X���e��n���"|H;!uL% /ߌ�} ώ��Hy��}� 0��Tb���G�gp�;�pCݟ��������FUrJ2K�j�LDG���r�N�2��1F@�dC��xH}�eyx�}_���'��3�F�V�?�F����-���6�|���L�ROS�DA�	^��6U�ݘ��ץ��rc�ݣ���i�Q��x�G���x�]6Ɨ�V����Q��et�Z�$��u���� ���ʲӋ<BJ�˿�2��И��f�B�W9�\��`a��`�C�Ջ'O!��u��h�i5Y�+����j�镳l�T�#�����z����C�'�)X���٪l���ԂP��EHj�݉�q���J��p;DS>+��6\�R��0�^R�^Q	Q�kЊj�j:&Q6,K�|�]8�xe����*SΒ�,y�U���P1n|@V���������#��!�d���[��p	A=zod������pDjڜ�0���L�8	_L��|,�!e����dAt��#��Ff P��"8��	��S����S�� �{������7I�d�n}��M�LO��ҦNb����O%�"S�O�&��F�T�y���ZN_�:0�ӡQ�^�A���3aN��v�0�������X!��x�&�T�7o"�J�eV���E���V��4z�.�R�u1���J��L�$�x8�1����ol�[�փ��UpƲZu�[�Pn�w�TG~ݏ��FT��:\�����[#�L)t7��+r�V��ԝ��R���zmJ���a�jn[�C���SK_O� ���5w�D)���r�|֊�7�b;fg�u5̤{Ñq�߫A�Ӿzh�ӏA6����͉Jl�󇵬?�_�����^6�6�~�w�H9J�N�8ݍ��X��@��"n��?��)��sև*�U�0����QNڕ�������[S��H�/���7l�fP�:!����� �n���x�k��4��)��3H�����6���{�[�� ~�?z��b\�&�_/�^#��D>9t�nڬIoFR���u#zB��ט�b����6��ĵ�e��^���_�0�)6?LԽ�7������]�g0�j�	[W=�����q�uh8F����,:�ɻ�]�F��6�n�� D��ɑE:̄o#���{���멜"��:��i/]��IB]&7���: �$�s�
ė�':���MZ3���L��D���Y��ݞ��'3�)�4��m���0����� ���Y;T���E�3�Ζ"֋�#�aQ�lp��h~�:����њ�:}6�N72T<�<�ڄ*�}!����~�I( L%�^�c=ߨ��A�ǂ�wi=Y���{���ŁFf��x4�q&��z���������Y�Hu}�G�
>h�� ������Tp�����B�f��ě�wb�kw8�K$�
霄@�iڢ�e3�����S����&�.�>m���i���Au��!��/AS���) I�0��%���SAI-��>F>��DiB�ѵr��8�mT;
S�����V�@�]���^���@�ǧF��������:)1�m\H��;kq���5ogF�j�8U��;��W�k?8
�xw��AL�l
z��G�`*�u�\5��w+q�����k�h�d�^��eZJ��m��?�</\�$�w����5"k޳	�Fo~���X����]��vG��f��$��������LǇ��[.��wK�H�vL����@�kb(���]�,Z�>����G9�S+�eg_.a�t�7�=���q�J�"k�G*h�i �����2{4���96CZ󲟺�Pm:��Y��K��Ǚ�ܡ�|}�ڇ_^��Zǯ���զ5K��l�f��l��H,�,	�hJ�Ob@�n���[��H�/.D÷�B�5zY�{Yk���6��Eh��M8R�*d�:Ơr�ǩ�/�xerfۦ̓庺 ��[�د�Bʾ���#5���(��׽c5i���S�л��I^JnO�w��ߧ�+d�K`5�%瀼d�=&[yx)D��Ї3���L%�m=�]�F��@%�'�����m� Rj	%�h����w
D��6-���䨯��t��`�<���x0�SS�� �׶a�;���F�'X�!�բ(��Ie�W����w[���+�C��=߲���S`c櫑�1ll����b�[�	e*������K{�
	?"�U+7�����S�%Cf���qi�T�K�F�L9oUdLW _�=B��%Я��UiΜ��_s�Ὤ� r��3Hؒ[��h*ԣ{D�]����cW���a&5��"��k6xW�²�s��������t ��J���3���I��w��z��"[�:���x>���$�y���afRz���UH �2��+za��s���éD3�����QV���<ZD�a�n�l3:yV�5�B4Nkx�la�}�Ⱦy���f�b��Bu���p[)&K�9�?b���W��d@��-]�B�seF��ޥ/X���n������lP2X#2HW�l���o#mn�����g�piu!��+��R+`�++�y�ZÇ���#��fVy�|_��n�ϕ��F�H[3��l'��sQ:w�ĉ8��S��|��_a�ǰ0i`��5��'|�L	�Yb?*��-����-͙7�q�L�HC9��+WWpq� �vφ�dOxY:�6�����T�� �|\�TM���(�vx�X���s5�/��M��.��5O�hP;�dq�<��-;+�O��DPϟ�I��*^����!Z�����|��5�F}��~�+��uЙ�G��+����B�Hi��{J�	�b�3�v�|�[oG~�xԜ�����
��5/W/�П+�$�k�5��k�n�qK���Fd�#��A�_SW�Kf�I�����(<0ޯ������ �l�����T	�_�osN��\h.DJ��]���:\���$�:عY=#_�^��+�	�#��BS.����B� *Q��(2I��wB�!��C"��\ȡ�xs�ܚ�Lh��X',�-�����.D��ۉ~U������.)4w?~Y�_oK!:���?�l?�+e�w�}3;���s;:��|��a\��3�z��@��i!�lϲ企 WzT�� P�lѮ�z��4�SN�+����`�GV�JY��9���V���~�K�[�떟�aG���_�zʿ�	�f�.~�`���<Sٽݛ�f�,$�r�Ŏ���E��aɬ�3���U�I�NS��OΈ�:��(;]�� �T4�G{;�k�������5��m|k��zURb(l����T3�!m��x<	�(��:�P�_����]��?D�!����||��*O[21.T�+�A�B��TA�����]� �C�����J�+��۽Zg���9�o�9&�3�Ӡ_��媜P9�06jxY����Qs�i4DktM�q���p���a���Dwv8(N#�җ�����tY���t�򍃔�^�\C�V�S�=a�$٨ĆH��W0j,:�`��l��O�ky��o�~0�HT-�5�/x+{��'.
�pW�(�}��bM�sQ̫Z����1c#"��瞥Sm4�ѵ�.	^�:�B��l�Jz3}F�DS�&��q�8)�<l�D����
��VYe�ǟ��^���m��gk��.֋�y�em�����m{�a|���,-���ua焨�dm�3s��"���'�5�@?t�7�W���Nݛ�p��i�rė�3�I�N2C��K�[4���f!5dS�s�����tq�{oc�աYJ\A�s�|��?���$����rϬp�� ����r�a9�W�}[�潐-�F�wE�;�c�li��L��	���$�T��4uL����/�t�6�pҠ"L,�d)k�#���3Xf�eY��<�)�,��Z3�Ȩ#���F?��ȞƟ���o0y�ܧ���F��e[�
GD߅� }L�~ҎL~��vCU�ۣ}ゔV9l��D�������-����=�h���ץ��d�<!B|-n �x'^��'h�ڷVQ�����!"}c*��a������婄�+�UX|� M�^�;���r��v����}�W�;��b���K��N�b9��1<I�����+6T�/�A��j���Wq,��!�tM�)�,x(C3u#uB����%5�+4d?}���z#ϻhNZ�ڢ�%�b� �������J�����]�V����b�-�۽�����˽i����Q=+�&%֧ˌ?Q�@-��i�/�H�����ҵ���l�r�Uz�TQk����X�WO�c�����������$���_<�p�2-o���z��D��Q�f�+^��X��ۻ���Dӹ�I�N��a�/��U����6lN5�������s@�O����nuQ=���D�UL���=]���x�J�óEv���Ƅc�c�Ӽ 2ʈQDd��ةe�30LO|u�Qw��$�S�W����@W��]�>�jʰ|��������\8��XF9o�5��>�(PĹ�X�~����C�H�-�]dD_�ϙg�oO��ꎫ�5{�#�ӄ�!��,��I�A2$���]�.�f��%#��3�f�r�����'�Xf�����]�23�S��R{��n���ٷ0�@�mt4]�^2��4�ߚa��Q�Z��e��(�H��a��'Q���7�+<�}���g�n�4Ju�n���|�9����4P6g�u�����K�\������A��7�e�R?��kv]`�K����Qo�$<D�������0��.�(���2N�������i�@��S�dwr�����P���:������:�7�3�47��z��pNK	-a*e$�����_�i0*�]�'d]���T59��-�e=�YrF�T C�+j�pD�;ܵ�{��č�[[���F������ᗋg�w^�%�J9��Fc4A8F;zб���@B�58��_�gJvm,�Q��1�%˖ -N�}����y�Ӛ�C.Mt-tx>b@h�_��ƛ+�;,V[5~��$R������O�Y�I��	�8?���@`����9��ӿ�F�~mQ�����'n�n�ͼeN�bB���'������<�΄�^��s9��DNQ:�IWJS���-��NJ+�fl���2P��F��Y�ö���\���[ex�l&mk������JN�]=p=UV�tj�6���F�5�t��sd�Z6��XΎj�"m�~���bUq�9\c��cNCZ����j�����!�#K�9���{�Q�_��
R B��F���Co����ٔ��I�χ�>�j�`�x��޲�G7��.}{A&E�ؾT�Þ7�dEJ���2}����q�� �?���7�
 U�fңr���i��,�~�i͝q���L]F" �xm����������\m�ľ�N[��ޮ�o	�Uyז��1K�.���Z�'��P1����hJN/;���s1W���W��o�S��$kc�\�f�9(�/P�W��Zd����nf���L��?	�mr@�$�ۭs�G�������i}���VҚ_�Ɗ4P���&��#�&����a^�E�Ux��<���u���Y��sN3#Ƽ#�a��i�؆E����&��Q�୾��.⋕����Ub��NV���Z��ńDpn�<ͣ�È7�&�g1�e��~	��>�����hoIx��L^x��@�N��Z(���O��A�bOd��/:_�������XJKbq�z�!d���{����:D'���e'���?g�K��ʾq��<� �����?v��gY 2�w4�]�@;�����=�]~�j�L�I�����q1�����p=�ǃ����:�(L� �Ǌɮ.�o�-���"�(�n�؂D�����"\cįD�?�(����%��|J�W�y�&�����*|��u�h�2[Ϛ��~i����
�N7�����sޕ��{c�q��xH�<W�>*Ux�4+�S��a���i�S��}�/���O��!���o��"��.��r�����U@���N߭!U��H('�,�j��t��+�n�y�K^�7�b-4ӆh�Y"���\ĳI�H��	J��4��̳Fڷɣѭ2�?�{�1�>�hED�9�;l�?�~�ه\Β=}�3��:,��Đ���j��<�d���8[֯�Fǒ����{U�i2G+W(���2��8{J��[}�Ol���|ᖻ�7"�z�:z%����9�f�A��X���Kl)�}���T���%�F���"��n�a��_� q�i��W!��1��麚��P̘��9��F��̤12�R9�z�Rz>Wt�f+�ò%
��@W������,�N�
�ys�6p��״/Q��ʼ�#Uλ�R��Ԃl����NMo�u��Vj���b�[?kO� N�<*��k�x���c��fai��Ͷ�C;���A�ʏ�W���Dp���(V�0��6E�4ႌJG�ep�� ���w�0�_�}�|��"RU �_E��KĔ"� �ȵ���b���ޱY�=�S=!!�����o#]�J�Ҫr�w�\1A�Wy4�wH�O������/;7$|�Ժ�:�񦮟���c��#�>�2�r�*� ��7�^�tYW�h������gR>�Z�`¤�ʅ��7ٱxgP�*$9���7�Rl�"k�?F��ʲ�ʨE��i�i�GzK�΁���0='�]nf=�0Z�����b`=�9�+u�ҁ��m4rFS��<��ŷ$Þ���b��&�kf,G�P��63����7�?�he��p�^:�:Á��,��
圄 R��6���z9%��A���P;���@��'��@��n��q��C��hI�M��mN�w���1���T�W���D�KX�d
���V>���ۭLe+�� ?�[J:D��b�Ai���:��D�1X7�>�6���k�o�?Z��/{q����^�[^hUӐ;� a�\�_��;D��~?���8+�f��j���/�� ϐN2ߥ�F�h�H���LHd��v�2*�߂.�f��ߜگ�n1҆�d�%�~����%_�����`��kdNM�T������`cYZ؇e��O��W��w��ъ��do�K�~YR>�����u>A����>�K��N�K��Qe  ����i���^'�Hq��*���T3�����ʝ��@�4�Z_a�Z���Ʌ@��k�fc.�Y7��O_Z�E�M�C�i#��渽`Z(@2��5���w�A�L���$��� ��9����vDK�W��`��,�H�x�����U���i��_�r쩥��T�SpP�!�k�*�6��w$�/�Ȉ��:��~6 27�v�S�����h�)�lZeQM�8O�kLD3�䏹���|L�u?��.�pD�Jk��U����Gl�/����ǲ�͖^Y]�_�6̄��&�SK������s���9T������E}�־0K|l"h�:Rf�q6Vy��"�}�u�\=
��!�HV�ޣe 76ܡ�] ����d��d�p��|���:�>cx	���U�,3e|`��0zlB�eD,PG֠�Z���e�Z:�I�}%X>�Jw�{;�v��X@ Q����+g/�D�x�����.i��|�gx&S�G�����D��������V�ױcv�ܵ4Z/eĆ6��q2�:1���(w�_�� /����.wd=9��/-���.�A�����	{M�}
��r3y��n���h��s�����%�T��9�"�|@�A?�.oS����>�:G�F=���{�Lԏ��j�H���܁��8��P8���! ��8'|Gu�)���e��wBL" �\�e#�̅������/��O�Μ��=��y�<�l쓧��B�)�tƗ��Zg~�"jӫ�s�˽��u.�&��YTx��|Y��@&����:!��=�o�o���#Ȕ��$��U��Fմ���&�}���.�?�)KKuTsV8 �گGJ<n"�5V�2�0�z.*��[��e3C���&�Yy�,m-�Y2�־���N�;���F�#���j�
q-L~}p��B5S�G��M��������םl�*xv6��T��2Js��^��$��w�o�q� �jo\B�f_E؟�k�/lj�����k=����Ph����ts���d�N�7Z,D����[n.a誇�E�$�4&���l=_�TR���r�����;L#����I��<`Д���!��k�r����Z�f���{��������sX��}��y|]����Ԓ̯����N`�B� ��A�
��J�^[��<:��W�-w`�ʣQ����B��e�l��]z��Ք�(d��5�>�RI�H}�5������Rg}��tQY5��]d�I���L��·�{w��MX�G�����cpO�l��r��6���D?>Ԕ�����H'C�`ޠ�G�o��j��J"n�3c�������zV�5�OfK�eǆ���B�0�3�&�������w}h�N�+oDD�db�۬�*�iu���#�UG�ʤ
�-Dk�F|����?�keY"�L=��11W[�Ԧ��a�[@����W*�����"�6!�fp2=c���L�g�P�h�\-=�f�B��<D�4oH����B��QC��ug/���Kݜ�9�һ�㬺�]�L^4�|n~�f]�j��WS/����+���m����.�������!����������Cp���]�}���9=էj諾{�hH���uq�&�y���󤪎��"�uvĎ�g�FC�<�n�M��ѧ��G�ץ��. j�_>�A�����Vk�3_�d' �R|����7���M9�'�������	��8������k���� +����$TX8*�.Rx��r���MI>�II�"�4�E�g�!�!&��;Z�F��ߖ]SW񤑵�S�ܼ��/�CA�v��#���.0Ɖ�q��M
�Dr�*������zb￙k�W���]@�ޚ ��8,��_S_��]NCK�F�Xw�۲j�[���i1�C��T�諾'��b�B_�.��.����a��q���?���v�E%���HA���`����h���E�/K�f��\���2�Qj���N
�'��cZz��UW5����l���wg�ɑ���@R��^-��'�d�g��
3��
(= �3�&�ˮ���|��^�9BG�;_&�B�y�[el�z�����&(��*�~}��p���љe�/o^*�/T:�����짚�/���l��z<���Ma�����`����w�����0)�#�[��� R�����:��5t��C��.ߢSȷVV��|���j-�T8^~Ne�^_���a}�� �d<0�N�AAv�|\5�����=>��|H
0ų ^�T��5���ՏD��r��|/'gĀb�?vwU��;[���_���6��/Oq��,�À�u\�`H�#�Y�8V���eؘn���C��S�_�����X+����w!֡�G��y�+}����r��|O�1:�4�7I��:If4AY8x@�|5�c��= (l���f|a����3�^�ޏV�5j�L`��v=xq�o]��p���s��NX���Έ�ԟ�$��a5����Xvj��G�ǏM����Lh00�!�`���D`>R�R�}��י���{Z:4_`�b��R!�_�U��.����P��G���X��o���@�SV�E.���|����?�C���qڧ��㭯XB��'�D��L�b�Hx�iĆ`(@�0�$�%q�J퀠*Pߠ���D�Ð9��֠�����yO�,=��R���c���0kmV|�^�w4��Q�$����C���Q���5/\�(�&	,Ƌ�y�1A�� �P�ҩ	0�b6z�T��Î4���h99����IQ�U��D��2���/��D�2��N�N|�|:+���O�A�*IS#@ּ����O�gS[mdش֍���~^���Tgt�)9&�G���'����R>dh��m���{V�����S������C���<��L$#)��#����>��������W�JHgk��]�E�2)��xm�|�/C�w�F�c�Z�?"�eQ #r��@���_�l�P�?���J}l���i6�ղL[�Yk0��5�?dtJ��o�H
�f�هܨ;�mI����A��bj���'�����V|ۄ�/ �!������E�#$�P��&#;� ��ZOO4�$F��>�e+�wT�m�L�a7Ne�����_�Y9U����	�Qُ��t$���g
2L	���T~����O�b�$��{��C4i;L�>k�x��F>�ێ]����ҵ�n�G��tS����m��7�hm��y����-00�������5��	p�z���cx<�H���f�s6?W�I����KG�t�0�|��+�5�N!����)���,�$n��Q�S�K�>W#^e�����k���=��c�-�����<f���|�U�1��ReV�*���ߋ\�ػN��`N�ñN��Q@�$-�2��+�$����L��c�n|R���g,��W0r�A2�v�����V�����W|��Ҷ#��㗬����{sc��1��|jd~�w��Ki�&LF�ZO��:c,$v<!M�b���~��?/c8��jQ^�Q�FE�>�������N���7>V��y�����V ��t���ǝ'po>��o1]c��r}�@��MV#LH�ʲ�͛��j�>���B�X ��Z��-�_Ӽ�_��h�r��ϵ�+�iц1ƈ-#�N+;h�"!�($k��/�5{<�3�[^^��
�4D�M]�ڄ������ky?DMꈅM|��-X6{
��~��N�t���
����A���]����bq��y��_��d�v��q_w0�~؇~�;���a:v���࢜�����q�L��sRt�.Xh���x����j�6�XIe3È��y{�C�i�3���-��o.�	��]6�%bІ�����~�t�Ѹ�h�7l��'�ʞr�C�⤣��i����ĊN�7I�A:pK���X���Q�5����ݲNf�)�E]�`?�tLk��WQ*Ӎ�Uؙ��vF��Q؀��n�Y�%�������U�q�N��4%q���}����o��F�����J=���V����s��L<Av��AbNhB����[�}�A?�-Re���<����(c���Ҿ�?��.��"��X+�1�mQ��B���T޾��:K�c�d�g�0��9�:�E��D�M�y�u��*U��CL֕K�v�-�<��m�_{�p,�JL�E���_�(�X�>3*K�p��aא9�_|�k ���Q��q�M�b�˴q&�2dz���q&;�A1��P��c�U���nU��M��_
_�u�B�}�6^�x�u�Ry0.�<���h� �����
'Y�ڂH�)��$龠d�f�ǿe�a�x�}���~���8#`��Z0�/���q����ёR���%g�n�''���@� >�K;���-���La��xA�/�t��T��<����)�->�9��%���s�˝��:�x��b@&�g�r��I����7��~l��ϐ;����Ư�:v�!���m�v�A�P�a��_~X�(�]B��@�Z�NsC�4���=�bS7�
��I~L4��Ida��k�.�>�cm��n��z,G9�р|aJJ6pn�O0�|R�^ؽ<mw��#���,SO�HK����#�d{\4��B������,Ѐp�LD�����o�;\�I@�;o�<�5���9�ɭ���ϸY�,}���F��qvHg��f5x�e˨�u�A��cA0t獝�%��λ���e���C=�t7���F�)�z���&�O߽��31� �zm75��-q���R��<�)��7��i�F�)�6C�T�CۼH�G>��ld�'��gG�~�`��=��Ms��Kv��t�Wq��m��q�v�|�WC<|2��~FcC��	aFX�w�1����O²:�`A�Ut�}r�j�z'7��GY��CƜ/���D�e��ZBu������ދ2~��.2UÜ5����&�1-ƞ���s�!W��Dҏء�V]](L����~e��c�*5�7R��_iO����az�����Ń0l���eW��Q��p�D_�F�D��rٓ�!Cy��2�)0�Mp��`޺s�죝*����2;p}c.�)>	��̷�dȮ�-�U�|^S
4әJ������z����t����)�eN2X���|��sPָ��
@�$��R��W��Wo��{+훊�����2�a%��a��bL�$!4[�i�?�Y�[��,����u)�ܓ1h^���BL�&R���>;���S�C�&����Ps�>x`,��W}������������i���A;���E��sC�pu�m��fi7��Qθ�C��1֠�m?*�-D%#�!%NaE�q��HT,f�et&�il��Uj�j�D���t�p|�RW�>t.)k"�r��BC�$,�BZ��/��Ct�A�}����PN�?���O��WǑ\��~T�������J;>+:9n��y� SpAx~�R ��F�|�t0�)�:~&K�A0R&=̤�$<�楖���L~K��p::�M������mu�ܹ4�8�r;�$�GE>��V���-�LPq��<��pv������	�ͮ%;��^JE��Z�u,D�Y����0���m�FS�2UB.Nq��ݑ��/����ZQ��h��C�}��:�G�HM9E���L���J��m:�k����L�M� ����\K�ʎy����P�Q��_��] �<��$\+#,`�9-PM�S���ޏV���K>�z�/��Y�ѷ��4��Tn�
�t0��<��9-t*d�#A{ҽm�F�o�\L	\F�!ֆH���	�-ן�G�A���%yC��]��V ��qɢ!��&�����XhM�%È�ё�Ϗ����ӣš�SfAN��F)M����	h��� ����@O��3b!����9S�����v�l�a��3N���r�o�jQ�`�6h����.6�R�_�I!��RI뱦t�����Ȭy.ZZ�"]��I�[6�AP�l�Ȉ�K�[*�v��/|��Ȝr�H��æi��! &6"�ZTKvo��6���L�J��ټT��?��~�| �f&�C�itn�D�=r)�g���l�~���͟1��P2D��<�$����o34�kAܴb��įU�vJ�¦��{ę�d�zw�z������m�co�&������B')�!: �h&���%�D��e��Y��n���J�eoI��aD���rE��fZ1���3�'�����c��C>i��6]�>N�D���fٷw�I���N����(��Ws| �d�h8��Ѫ���Le^+]��(�q�Ό���������du��@��*���W��=�稱d�1�j���5����Hci�x�O��r���Q�Zt6�=�oUZ�P�?�}׍r���3�!P˺Y1�5˖mYg��XI�CXi۰�+�,}�"�h
��o>�|3J@���N��'����f�y�g6p���J�����j]ꤦʂ=�.,U�e*��Ŧ���VqO[�V���Ŷ�v��O#S11oC96�\�z���8�aW��#8*�5���LCj�}Idn܆��1XI�_x��������2�^�<E���٘��d=���&��"5��"��� �2M��i��	���\�E��DDG�OVs�,��N�<������,c	�±��V��<@
��~���7E�gom��IS!;y�h�kd� ��^�&P�Gĵ������&�.#�|�j'mw>=\��H �q�X?&�v��u�j��R
�*߿�v}�h�d��Ag�ވ|f����U���-�2�B�g�mY
�xY�����l��==�p���a��9K��z��
`��4�Y�BN�Y�3m˺O�yr� 4�v�o;�F�ݺ�=���7T�(=E��V?���w.�y��Y�C�NrXh�G�<{��}�#��.h�3q�-RAw�\�s�ϸ9�!.u�[�z��T<̸q2�ú�HH��9�07���Mi����v��0���G�Q�`�J����������#	GsA�;�B{��ƭ������빱��~0\��'�p~��O�o|b�|��	GA�Rooo�h-�k��^[�N�?���-Swj���m�q�k�N'�:�L���~�Z9�T��g�>З �0&Ҋl`��}���Լ���f���(%�R����Z����5{�ſ��?Ӿ�y�����([T<�t����y�o@I�-��\6Y�ݼ�e�e�zv�)��g#6a�Mt�M����D�Bp��������\�O�b��P5�B_�n#;��8�@/S�y �F@�l��}|t�. ����k[	�:� 5�J�S+���8�c/�Gl̂�:bt��RE5O�.��h>��ײ%J��z�^�%Qr�����f5�Rt�8R1F�`��J�$~3�edhG)4A*���B�I���x0��J������r�n�)p-C;�2eP��� ���5p�2�Q�6)f�,��!���+َ�m"��[sd���E�o2��=e��u���^�V�=	ߘ[��m��52-iSx*�˳���ӈ�\}?T�f�����-&(�[y (����c��'n���pڎr��n��f`]&cO!撲%����NR����:/=�%l�)Ȇ��Oh� �|cS�K!��I�b!�|L��XOX�׋�H���-�6�o\ߏ�^�B�Z���N���VX��CVn��GgVy5�?J)I�S�� h%x>R��NM��Xl�џ�;ʟd�:�'��t��m�F6���}�j��^����o���A�ܷn-)�� W�$;? 	��(�����U{*���	Hx,����G2e�H^E��Z	����g�v��i��t��& I-�a7��$=��`�G'�7�\Ym�	2x3�x�V�[��J1$!<!�e��r5�v@���[[89�Йl�S��·/�ͯ��Rݝ��T��1�30�|�:�Y��*	�����"�|.��Hd��W&n�gLc�#����W�K˼�/�F�f0��uthO��糰��<��ya}����M�*�EPM�z6w��s��ϮZK�͆�+ۄ���6	�xa ��D+c��1�eF.�-$���t�fԁ��$����:i�u��;K����.��3��M�%eWlu=�Ee9OϞ�!} �H�K3���5��^I�� AGŊ��8����E��@�M�{`3U֛m�>e�/���bU����,���}��₎��R*����=d��V�`Qu�?�e����g��� �Ӊ�&��QP�ibI���3R�j����4*��T�k'��I��cezǩ;3�]��7�p?A#|$�\��o���J�����k�5�#g/��j�>���v�(b���q��$ō��V�	�2��wh�f+N��k�f���
��w�����N�_:�z��Sq���Ez`@�#u���~�0�SQ�'���E�����N��[kׇ�!iJC����J�-��7z�%g<fJ:���|:���ks���S������?G�j0)�kc��H�#8{��-���BIߘ��̿��������{k2#�v�&}�]ca:�-iF�8~�~������������}�Q����묊�OxWL�Ð�i�4��xI'�yw������I����z��J�۪��M�|�uނ���&� 2N�(�?��mף0�����)������kQ@�T?�fU���M��2�S���Lr�D��8J�"t�!s-���|eĖ�hZ)%x6�(ub��0���h�c�XE�x������e�5�У�4��0�*�W�x�֪G��]W�3W���t�Xsd�t�6*�����W��j✅:H����{��펀Z����d̭ω=H%�N�'���{�B�{}�RJ�yxe��E�\��t�>F�bwި�꤂;7�/��(��`5��A\��Y�:���	_�&<��qp��X�u�����ǻ�W��2d1
��'�CU�5�ۥ�ا�X�,�����R �ns������sԹy��3��i�����.4�p�Z�V�K���N�2��#���W7n�v�}>0L9�}�SV���֦�X�.$��8��jM0O�C�-�l�*V�6��uӡ6����	�Q����o�C,�LZq��b#�2&:�?��`^�vS.��`q���B``��8D�(�˄�	p��8���&6�)`vA���P2Ui<��ܛ�~��P��ݱ�#����|5tw*�$�N���L9���˒�lg�]N9��!K��Y}]o�Q�z3�F�N���fS��hZ�]�8��ï� Ş̠����~���T	����x�l_#=�ʭ���ѫ����%�������#�Vv�˸�ĸ�C��K���@�J�h�詤��E޽��-��S�����5F<���2 2�������o�x���y��Y.h�ݙ�*���2s2o���Ȉ��8���{��C [{ h�M6c	�!m`m��bs�����`��L̬��u�t!�`���>�3Kf�d�93!*�5����|�W��*�CB&��3d�R6� �頶��$u��/s�.QGe��x4K�MQ6�b3����"_	@��c+��]���9e3��4x�`��Uo-����R�w
G߹ʲ����,���x�Y��^g�=$+�V/�1�Re��/d����S�W/_��D����[�?�	�G;�"�1`?���Kc���O�z(�Q��]��&;��4��hJv�~Od	m�DJy��uL)��-©������n t��"�������|s5�3e�1U�<#d~���N�#��!y�&&���#�J����G{k���X��ǹ�(��D�ɶ�4J��r���O?���`ا�@*�(�� ��o>o��|���,�Yg������Ig�\eɂ�:b�0����P^^U6֚/
�!��D�TO��j%�K+��h�on?�/���2�nkݵ�9u��o�8ËE���_H�P����2yM~֐�+S	�bq
GV^{���|��s���-y���/-��bX���	�t~����j8���ؽ0k���M��RY�q����~���.����ҽL��U����/Ť���o�}�\*Ǭ͡�0:\t��Szj�pTO���y��¢�3��al@!Fw D�J�I�̓�%�ŭ���R��]�"]�@�y@QKaR h�R׃8)R �'���"[��[���p���嚊��
*�(W��_���S��HZ|������#n�(�ܞ�6X�V�%�ğ:���-�]t)­�@4����&}��{nE��2ĝV��JՎ��t]q&��S�\zL� �����C�(�\N��~�j�8��Ř�7%+a��ܾ��m5�e���X�oA�5��3��_���Q�`��=,Gez�4�_o>�<ݢ��\��9GV��YXʰ[�������`X�f6H�57�w�+��.��a���{]s��2xy���y�����wgD�M�%t�rn��"e/���[�g"�?[�	�Go����a.�J1,J>D�:��g�F�A�ι��87�q����s�ñ��f�Hz]b���@�-�צ�cM�Z?�0�Fv�	��@vҸgJKkBm�%I�.���a�*cm xtM����
�#�,:(�oA4����6�����a�{5��1nuuxJ����}Z�j��c@t��������OO��(�d)�e_v2��UJ�q�2�{t�ɸ �˓|����89���I�KJ��=���c������+�fāݩn���lO���Z|�D�il��T�c�: i��y頿���t���L;=Kur���j���/���w��F#�NA��'����<#v�\H�
9cӇB�i#EVF.���4�mN��魩f]+����� S=���޽�O��1iI�����������<�������h�wh0�JB%V	�7�w��Ƙ�(	��Ղ����;�Cf;o)�����F�����0��dB\�Q��������
�_����r_��[{>�Cꔵ��W�9\�eT�u=Ʇ����3q�R&Z� �A� ?����3�E�х5'��Y��5�r۫ɚcd��<+8�Lo���X��d�q��@qj>/�X˼�pÆ.�i޾��RTN���wz�n�����Y��\N�`})��d4��1��u"�����5���XDбme|��a��{��Y� �7-�~�
X�uc����ѹ ���Y�B�|k�1㥔�iV��V[�J/D�ө&?{{<8}&�n��ZV�̜���:a�U�a#��)j�
�wi��u���a	�ߛS��}�$�c^3����Z;�Y9���'>�F�\�V�S@�eί5���Ȭ�r|����NV=S1�� ck����_��S� }�Wз $�x�ij/����q�K.�Hր�Ia��x�^9�T��X)�����0	�����������f��]��A4��*�#��C�˭}�mz`���N��O��A��,۟"gǉ�V6��2M�va�ez{��?8uyJ�[[y=
2�C�e8'���n��\m�]�u\sJ,��l��C�s����`l��e]x�ަi�?�	ӹ��5j �"dr������5cQ���0��M&���N�$��OiZ��)��C��-l2�J����T���_���\�2��2P��R���ĺ>�Gxv����DS>��m +��R�n=A�^�ݲn�(oi��>�͈�CWM^�,�h�߂x�d(�y�?����D_��>1�ɱϡt�����d�����H T�Gַ�M�A��Ӆ�oF��6⣩&A����Վf"=�����Y#l�J��dn>��vR�p����f�2e�0Iwl5Z4�7�\ �7�|sG:�b�΢�R��#�[�6+�AZ�d��'�F	e¾f���*K����/���Z�RѮE�~B�T���Q�k_z�g���3��=L�j6��et�Q�I5��#�kY�^�Թ���Kzy�#ߌ$�*�}T�a����ڏXi������� sl���C�:��(<Vx=JՏzuĨ�3��V���Y�S���Q���2 �#�\�A��f��kK� �p�������%�8� U=�Ξ�i���1��:�a;���;у:H��$�V��YD��ҷ'�J'�A�Vj�~�"n����DP��Ғ�m��VV:�����>�j�Ҡ����@�>��/!���1�sZ�6!�a���G���x|�jh�AJ�i�s��yd附��!`���J\~�ţ�#�v�.%�5��NM'�3���F�*j�|����H\�[�gs���cO1g9���D'F���=��F!�g��U�,mi�ώ|��v#x�5\tM��ݿ�5�Dd�u�_{ړWr��}������k��[��-�	p�GB�D�eZAI�V;�rjA���e�G�ȑ����i�c�u��\�c�~���9��pP�J������� �amvC��-j� cp�Tl�x����먡hΟo�����uٶU�4:�:��3C#"(## �i�J�Xa����WR��D){�X��E��������tYy�9�w����X����ɘ�1g �O��7�xX%=����p+�\�d����hi���+�Z���b}5�ƍ�[D'rGx6#���b��N�RP���S�����tW`5�<�I�h�˻ɟ#_��F߾ֻ���C�����th�߳�F	��� V�*��_�B�����{��U� �\�v,&�۹}�z�_����%�Y��oj�U��p�k����x�k��clғj���2�_����J_߾�r�~y��'3C_��|u��JoH��^��\��P��3�:4��UO/I��jٛ&�I���Y�1�Y�/����7Oq�c>wQu�H��){aB������&�jOg��b������p����ݷ~�l>y�)H���$~�Ž#;\�	�.�sH��T]�G�ϵ���G�u�=��=ew	J�[d�c�z�fF���-�(5¨A��]|f�z�*��Vs��H
����Q�NL�o���'�?i>���ۜ_ȋ2��+Z6��]o��_ս���ǎ(8 ���P(F-�i��:��y?ߞ����Ų?��$O�E?�� 
t=U3]�^�K�S����,OF�# ����c/ئ+n`�fױc?��<_�7��xfn{�}G�:S���
,���|�P��M��Tѱ�3��1+Q�����o��5�z0�����<^s�Β�����*���N�IlY��zNd���v�Dl����91b��-�Փ�bEڞ�����#�4��'n�2��Vc��[`�ZcF�����DP�om��O��D�s��*w���-p-dS�Б��t
V���5�n:k�kY�W���TG툹*J�(�m�/)�R�	��|�bn����/ۖ#��&Q���P�\���>��dMeU�/3"�6�p/���L�|�Ϗ�X[���Vʡ\>�Apd��W�K�|7����6����Ӗt�a%�Sn���I��]#΂����819�I����*���p+K���Ů�6���1k��Pp��6��ی6�w���B dl}���F_�h��Z?8�uw1�S2ב�d6������t��:����6�� �ˎQ�����쐮`��ps���
׮z(��S�#�+.��+\�j�R~�����>����56�Ҧ�\iكPS���$Mm9�Qb4�F�o���e���
���zf�̫�yː{�R8x{�����5��Xu�O�U-�վ����b��1�157�=�)���Ki�T{���~RC]"�h�J��Lc��z&wz_bĴ�UG����E��Q6+n�m)�-�iwk��{c�[W�5����#��(�	@�ۑ@������(�J�;&��Ңe)���I���xA��Y���&��i�^=� ���5|*W�WV�JTpk�YgG�XmgB��`�@�E��lk���t.��9	���^+S��Է�\���lY�	�k(��M5�i����zٰ�о1�Έ��uc����pyK�iN-u��S(0l�w��P�	J��?C3�e��6+�ٕ�B�՟ �.$V�C�	��'oF��}n�6���A� ��G@.f���U64�����[��N�c�9eR �
�~B���a�#�V�Hֽ��Ҝc ����y�^�_��~��`��:]/���l�s��˭��4�v���*|p �DX���8abe���7̭���ܳ�M�U OvVc�5�<O�w�x�*��(H�|��c-)˄o�>����]�'2_�?}f�a�&���46O�&:1Wx��=�12��{��f�lQi�s���n�#�U�{��ʋ��7k?#�4����9����R���pAj�r�1�ˍ�b
�i�������n���!���cj&�|;�D�ʱ��+=�A B
oEӧ�8�*������r��_�EF`}��[���F"o�3�)BJEKS�6;ΰIp��8[���E���U���(i�ͮ����v�i،�CC%������u���s80�	��������)=w*��͂��Y���!�6�Sj�L�I����4)M�H��t�%�d��F�ɚ� ȱ�TH�J;��x|��Oy�ش#���'��	�jg�,�{���WӟUg�ȯ�^��Ts�q�t���B�+����vK��4�$��DC��^��p�oO9�b^�������s��}��k��Mu.��r����,�w�f)����l�2����P�줒�5�0�um?�AT
'ެWLO�?T�B �+�k{�&�!�Fu�a��*i�����zv:,y�͜�=AB�m�����ci��مɷ�Wn%����K��_��fI�wѰ�-���$T�*�mX$��7��+ɰa���ZJ�~;.���� ̓<�M�~�#��!]��[�l�BF|�3�%7'��@��iF{R�6�o��Ң�:h��գ���݃�̟U��ss�4�OBz.7өx�D����^��QR�#P!�E��k��fBmQ�ܛ��;�4l#z�u4#�q����%1<F���?�,��*�]�w���Y^y�zK�@����V��Vܫ&��UԘy�,��M�u� Z�(Z�SD'DF��h`6�bW����Q}��_p���a6�l�Fp��{t�ajHɸX}�Et�������}�x�Y������f��(�x�n�������gӴ*���>�w�ef�F.)����֘��/&�c�03����^%.�x��+(��q�i����R��Mӆ6��@��8�전�4��p��U?|�o�Pp���t�4\���-i[�%Np����0]�Dj����ߔ�7�v�|._���e<���}�x."�T�.An��H�a(����j��<bVz���GK�s�pS;7���E�fr�-�I�{�k�nv-²���ς]�O�|����)oռ��d�lU��d a��X��
��I��7�ג=`BxVn��|Z
�y�Q,Uo��H�ls�m�CŠ��G��Qx�����"��/�/h���W)R�d�5���BѶN��S«�QM�V�G���<��C��e[Xު��V򐓫&Fg��@w���S.�R�	�f]O�L�~�P�%:�7���Ϣ��	�hBj^���.D�\R�f�j��-���j��-��d+A�~��m]�LSaGl=��Pi�����e[�yo4�J��_�!nk޻���*��>�c6�rb���,�o09vH"c�_Q���m�&ܗPVL�~��k&!l/�b�r��p:�����Qڼ)t3q�U�O]�=Nr���!v�U���2�G�S�]-�B�\=����f�O�L����V~Ҕ&�;[$[�/le��&.Hw��3:���x�l���Wnt�K���2�\ׇ�.՛Z�/e�8߲#��������EMv:�)�^^C�{�$E��D���eM��d w�}Q�9+��S'�sh�=5��]��0m�i�X��{j��i���Q�����(c�;ߘ)��#�����m�VL
t&Np�mĠ�O�ǩO��2z-R�.��Y��6/�
O�v::���it6���M+��d�����۷���B8ꙢQ�6�C��C(	#h⵬�]
9�~[�	*/P4SrоC��>�A)��T��x9@�B�h��z)��s��t`E��\��?��Zcȟ%7q�zF��V�%���n���b*���$�0M����G4ח�nz�7S�Hy�ɡy��\;�6�^'C��_t�N���L>��TE�sZ�nL��-d��r��j=?��� Þ��A�_3���;�䂩���#:��Uލ>�l`^o-n�ܡ�:j���O�v��a�&���!-6�j1B� �J��"�@���#է��»3����������	|�$�5��U��ōy��
�x��qՎf�ǛJ�B����+mA��E�cci�����_Px7`���- t��/�}?C;��Ώ�dmT8lH�9Z�E��j�*
�n�6��5)�*"�m�5O�Q���3TZ�n�8V����/~�b��7|���N�e��'#�V]�&�v+w��U2�b�s~_��VH`q���O�x��n.u�������zHb�$�����}y��6?������h���\��[�#��S`�����#�=��i`�q�uS��+�Jv� �o�1t�6MR�4�Ac��m�;��wY�7��Y����P��o�ꧻ�^��=�4M�N�z~M����xFrGR􈦵�
ų�|�3 5;E�	�Â^9�(�:� �u��L�&�ck�hƿ�b��˔hB��P��A%xJ���4��9���p��JL�\^X����kW
�:��4��f}C����������#��,���u֜����^C9Qӣ,X��J ^���� �O����ζ�*����|�s���+�%�X�~�]mʜ��uIC̪JL.���ؗq+�!�O���n1��m��A��3���@S:���U={��Վ���}��P��d��y�6���+s_�zG�-���)/��lk��t�,����3�.���w08�9im�F��>�I�i�Y��+����>������A@⊵�F?=�X+�Ҿ&/bwl���5� ����E��e����M�M\ ʹ��Q�ԋ ��0��%OM'��inK�Aؙ���s��s����26�J�ކLΜ�(�/}3O��Q#J�Q���B� �D�����%���f�7̌pd�B���� M<�~����~�
G="����h����|3_��e!Λ2��ά��x�� ��o��,C�3�+-Gh���~�@�9a
�
�@���gI���"���ǯ��G��\^'8̊_�A;lӔ���3#>ϼ \xeiO3K��l����=G��8�� �	7Mې�C�nN���}�w�&wJz}��"��a��ۋş
���"���uK���^��֧~�aHޏ�~�-=���/�� aɹ�6��j#b�씩� ?�����%��tyvv�+ѣs��8̦��ٻ$������A�=ǹ���K�������Վ���/���;����k;
}�����`��[wq�@H�Ow�)��~��@˳�4�����/jH�:Y�(Y�,�����o��#�	w���iΒ�׽���;]��3���#���'3s��s�\�U��I����t�	n�(�>rĲ8ӽ'��iJ����.�Jy���d��X�`�m�̥�����X8��>�~�v�^���Ғ@����:��1�w3��5���li�k?����m'��[2-�+]s�{��俀�p���8��c]脳�����g�D�o���a�k1�"q%70`wd,eP`U��MHI�O�+�/��](���(|$��<��т�_�뮛]�>��zzp�=p"#���g�bBj;�+����-wI[} �
�����օb�/Fm�+�V)�*|����@ _��:C����RmYX��p�-�DB�7ʘux��`�jL:<X�����"�/��F����@n�M�#�cdU!����7W�}]ߘkb۶͉m�۶9�Ķm۶����߿�y����u��{���鮺Na��h
)E�H�֭cɋ8�~�6�i����R-o��i:�$w�{����M�oVg��^fv�P�:Gc
w4�~�Zi<^���\�q.R���v�$%ZJ�	�E6��~�|Ҏ�w�!1�8�:0���^-U�d�#��+���7�֫�S�vtQ"PB������{��N-�h�>�Ʃ�nwY/!c��¹��� ��d|ɉ�<�j5"�t���W��h��͑Wq�Ĵ��]ZG��^ye?�o ��K�=H���,9m{�q ��-�w���%4�1N�ϯ�ڭHcn�D�ܠ�t�b���*�vzk+���ԟ�O,�o(s=x��&�L�J%���NRʈW�d�:�ecU��\Ɖ�m䵂q��|��N҉-�̔��O'Э��OcR*^ǃ�5e��_���@m>����;�r�Ƴ�{��;�:[G��%��H�6m[�Ϡf���t�'�I��'��=�C�6�Fgd�x�WP�{�(Ȓ�����
u���
m���1X��]���@r�((��A�T������l���]H�����p�$�8"^���w���F�~�A�ִ1	�@T�	
�>�X��*n�%O�����c��d�$9c���ؕ��	#�B�9�_Å������Go0Y���'� ���p_:�}c4��u�.��5�b�'	�����܃�0�����am�<|�v��ɍk��$��r�0���?����C��͏>��5�&u���^қ�8��*�����NZjW�����Z�H�2�{�ԇ��Z=N������T�3R4���ÃX��i��ɻ�h]�Ti��QN�j��b	�%���t���	�\/��f%9>쨰Rc:�$�Q�������4Ĵ�Te�����/z��+�e�O���Ҹ��P̢�i�8%ޔ���p�5���*�|0Ҵ��,�M݃��Y���
���wf7 ȴء�!$F�'{>=�I���J���L:��&H�y����cK�#"��w�6����{�`}{(d�'�]�r�A��v�Z�i2�Dˤ[B|ͳ�����fP����淅���@+��V��̻0��d�&w7GϠ[�XYkTa�6��a�kPCa�0i���{�,a��ʬ����r������@f�!���� �#����1�_]���#e��9�Y2��X�B��N7�Pll��m3_K�M��<���4:��[������v���������c��EF�s5��;���/U�GZ?U)��g�뢨�*��1�6F͗�A���	7�|Ѯ`�)�蝨�����oś�1��/I2��Xv+���-D~��_Nz��'Ѣ��MC����q8��Uه<F+���a�n�[H��\�)%$h�X�����+��h��>&u/6��ç����'��W�MͩZH���ÌZi��la�Ic_ysri5�A�cگf�>��HF��{�>���` ��ໃ�Y���l�vgV$5[,��F���7)�D���{E�nh�2�O��0zUC>�����d��>8���l?�x�c����>Lh�5fhd�J��Ț��~�2m�����'��մ�1'�9�uԑ|�QXA�M,e�.�'O�İ��=��@�*��G
��/��:�7W���D�˷e���P���~��S�	���O"�<y�d�.Ng��K�z%>�	�;�M��o�D�M�u��ѡJk�?�9�G��l�ݫ��7�A{z��
��Z�j�ǌ��b�uo��X��5#�5�Й����m�>�8�R�����>�4j��Kd��`^���]�75	}�)���̌��
0rg��9�OB��%�Mw��)�k��+Z�ˇ��F��/�L�eD�z8������ k^�������;�\*p�5��|��
gw�|F�B�ȥ��,ћ
�U;O�8� #���dD��%߻�᫴�f�T-r"�E@�=������fi�)9*��#5&����+��\��Ч�i��>0�P!�Y����C|����U�'��w],�-s��F�����B���@��ہ�!Kۻ���&�y�r,��?	�G��r�G�2LF�N�hɒZTuӝ6t���U�$N��qOb�Ў��a�T{�/J��U
��1�yȄ�6��w���>"�f>w,�{m��[p� �}����Q*zi\PA�t]^�_��L�W�V�g��D���݉,�}�Ob������&�I� A����6�G��z?[(=B}q��.l$��U �q���~�`"��y�?�5Eȟ>�#oĕ�!���0Ɖ�F_�R���G|���DQ�}g1��G�ڗ�~MG���,UD�5o%�fWO�z�G�˽>5r�3H��OI����s�g]+�r���9Ȏ*}]���G�H�#i�@y��f������ae'"Q{��z^��L���iz?)�5�u�V;5|��]�h�z코,���&�=��|0�=p�G*\��P�̱'p \~G��������7:����i�3�t|焀���sh^�DJZ�X=�Y-	 ��jM��j�}�O�P������������(=�Bu��
��:om�}��r���)��3�/oOU^�������'�P��d:	��������WS$��M�{Y[���23>b��v��{u�S�w�5�LJ�6�:�����ﰇ.8=���'A���!���ϣ4	kԶw'\w
^�j��l 3�S���Kv����������5�� �GǅJ���H�����p*g�6Ґ����|s�R�DQ���
�F�11���~���q�F3�`i�!_{'N���@���{�������0Cr���.��t��$$�%*j�[�;y� _�����4۩Yٚ ���p5?�8y���A2��rS��_�<�6����K����?vd��*�z���;�t�(G.0��Ie��[�/���ގu�jb x+�T�`��lS��8�u��+�Ғ�ש�̒��)�X��}��=,��+�E?�{3���U���q��g��I����?]����a1sc�@�IA8Q"��ί���]�'ns���֥��^W/��2�\�4�;'�>ķ�	nn��0��ĭy�f�J5�B"¤w�.���w/��C?��)1�~y}�Q���޽a�g9��N z'������9)�� !S;Lk0ҁ���Vꁘ��7���O�O�bI�޽jN����9�`�]��ԟ�	p>O�S�&	�e{|6f������laNJ�#>�AF�gZ��
���R#
�˺�~a�Q+,kz!��UZE�gT�I��C�g���џV�z!�;wa�M�h�NDsx�kPi뻲�ջ��I6u��#E]�б�"I�r�!�zy���V�;�.zrO=���{:�X!BG��p�{@b�zǨFC����w��X����}|3"Y����|5:Ȗ�:O�:Y#�+V�"�n}����r���m�`����uN۩WŌ��� ���c�
k+���ʮZG�⽯�*���a��Čs�T3@Fq^W6yx���vR�4�`��#��<���i�}Z��.��c��>�}/~��ف��%�[���n�-BX`��<4�$�%�Gb�,f7��80޽~����g��n��X��r��"��zZ�+,(���ள}������B�/
�<�� �{X+I21�C�n&���G��3�Z���Zo|r�Z�?�e��t�l3&���Og�7d�Ĝi �aN�"r)�S�<����I����'�9@N����ER�2���y²��J�S�*^R	�f�������!���v��˒�ER����mrv�@A���+f�&	ܳ�
�����9_�i�8~k�E��-ka`Gy��t�8���^��ׯ	�l�
���Z�|
&�A�U>	��̺|xbr@M�2�v���AI_S_��i�|��d�|E\�^��$hI���ċ�048������!�<Z�4J��pY)Gt��%�� ;i����n�PǑ�?����Ȉ�-
$	����\�yR�����K���j��q�QP�$�1����ҫ�L_h��>������q��b2~w�9b�D�T�Hdm���tE�b>)����<�|&�@��o\�����6�"9K���p��O.06�[�J��$�i��Fu�Ң���Ko�p� �r0/�C&�a8M�O^&���������u �R�X�4��2��[l�^&>L>�%�Z��ad�=��L^Α_T&	+Hx��9�̜�Nv7cB�zl|�CR�&<�%%�h5=�|0�$��d��r0�N�yEe��ew���C��֩�� ��a�+�
C��7c.�mv��^�Y2'�������:N���9w��[��������re�����\)���o���!�a����\�t0v�`""_��DH�D�9M�U�P
��!=�g�W�LuB|��(��l��ӳ`����~%���<U�B�L��:c�ȧ�lN1��s�H���vR��ʌ��Q|�?(lt�ߗ�Sf�,�,wg���be��LMM;k6*��)�����f79u� i���?u�$�[��	�Y�"��K��L�?��]���c�A�\IL����]��:A5��c^�9�;��VKV�� ��w�֭4 �U[��E��b\	�3��2���,JP��2��d�p���_Z
@4s����#MM �N�H�83?uGYE�ȷA��I1kT ��0�a�O�����EMgK}5)�����'�}�Z���I6/~�Q��~F0��`TI��(*�C��t���a �SJk�����$�;}v�`;�7c��������wĶ���A���=�%rZ�,���AeS:�d���v�0<�2Lͯ�����:��pH"u�]/�{�*Ɔ�&1�"cL�M"np�M�;��~Ԅ���G�1����柌�q�~ΐ����b�T����]����i� ����̓���Ϫ*l~X�L�`�h d��O��_�X_5��˖:A��Lj�m�=���D�]�c5�6g*�rf�89�M@o��` ţ8���Q1�U1fg{]����O��qq�ٞ��\�:����b���~��H㺂�y&��KY��d��3�Ma�ʉh5{�K�p����@ÓUQ_�|U�,�)����͡��ͺ���8����W�w:p:FqJ�[�����}������=3�O��r�AP��3��Ŋ!��&���I�&�����)�C��D4R\6MX�2�߭X�?���.�< ��]���@@#�/�r*bĵXP � @� S0 �88���R���\��.z��5��z�s��	�nIJ';��_�~٩�!)P{a_��8 ���K6%���S'�w+ǙGt�i��j�,����1�i8�T�2NEuJ'��D���E*!���>��_~o;��|�uЪ���?�8z('��[���4f=���kúЇS\��%c���٬b6#;aB8���/�ޥ	�{ �6E��%.�lf����}����L��/�i/yD�E���-SGV��������v�2����!�/X]�=���L@Z���������Z�����Y�.��,%h�a��7ءb�=��Z�e���v��y�}M֖���W�?�����<?�5�Nc3i�.�0T���jɥH]��n`�1��㣔�U�� ��W�`�~`Tp|�q�@���fB�����ןcP�F���I�i�\�v�L�0ʖfMG���� �@��/p������O�.~m��)�������%}��L�s\_j��Ex���@2m�T}Fk�+�F�H�r�Q;xi�?�m�}�<�ҩ��o����Q�5N���d��Vt@�{W�:g����wL�3��_�6�L�N�+5�ᮦ����y�y�́-�[�Z��︧@ ��{�[���u.�	�0 N�����dq1��,B���$isq���mS!g3I�-NL96���Yf������ܢ��U �k�g��̞��Z����D�F�4�H�����wQ��o�vt@�\ZO�Y@GF����u{r#�hl=��Kf�M��]��J�̗��:!XJ��O(��	�{�6P]����=�C���P�V�([<;Ѷ)x�7{Y��|d,��0��9G]�4�FOO���IB ��s�T���dȐ��l���@�F�pX���:�������dF7u��ȝY�DN��ˑQD��]���D�k����r��pY����i��œP��o,C纐���ƹ2��I(b�W���,�߫Q���ʆH���=��~B���d��3E�$z�G���X�͘�$tj�P�T�hwU �p{���	���=Vur�� �;����cG$�"��mKϔ0Y'�s�䴏�p7���m�[�+�5S����G�q�y�����Ne������o�']T
m�j\�`�#,k�}�
^�$t�ڠ1�뙗������0Hx�2/�߷ '��� ��7��1T_��nش��S����㽖�VmH\T�V\��ȤpɈ�8�V�u�E>mrTcd|@D ۯ`�r���$m�M��^��Ձ�Q��s(�>�jO|�����&(w�?T��}Ƀ�K�|�/��*�- Pe^)aq>hq����O��!��{��R�ޞd�b5ݾ��ؼ���q�N�x"~�x���=0@j��B��(�t���m�?��V�`וX�W�'�A� d;���9�(�S��=��HM����&�}��5��Ŋ(V��Y`���`!(V�6�x*�d�{�λ@3z�n�7E9��� w�/ �#OL�'��B�oP�{}W����T��'��u�p��W`�@4k@���(}y�C&��'��&�����M6���x�l�K�9a��Q�TaD3&�F�7Q<7l4�B.���2X_'H�H���Z�i��2�?*;�wm�3�s�8�v��z4$80�3~T����-I:�"����Ns�q��J1>�bVd�������F��h� o˦i��kDB�T�zJ�{�[ �Le�t�a|��ɗ9��* \�k3S4�؜�N�Xzb2��Ȕ�;�Y��CE���z$E[86�;��͉-m\�i���Q{D$G�8���Wi�-�D۹R���ڤ����s��فi/�e��1耙#��#Y6�YJZ�A�ǌ*.�KM'o�K�X��6A"A
��%s��$o���A�'1��m�P��vgH�J����g<T�.�������F0�ug���c�����EAߊ���wG���-h��N��0�F�!%5^9�ۜ���;��#���sm�/4����y�l_Q��[���j���}R+k�|���)����o$/-%�G����3�2[<�>��i���;F����L-��)��[���938cL�S���"[��KA���=�ԟ�5Gk�{�b��Oj�;;X�/��\Y�DIl�]����B��_5E�M�'��Nq�I���z���rT��9�ֻ7��h
�h�)-fk�	�f�)�"w�յ�-.iEZ������"�Mn�9��FqbL��i�.�X��ِ��o%M���SQs�ͭi�'�m1�E�yŵ����]tR�*� 4b�-e�����_ENUD�f���D%���r4L���7}��$��?[��b'WӴ��e)Դ��^�q��Ѿ�"�y]�����l��U�ѹ�pLi�H�B��(.�͝�e~¯K�����9�C�V�_��Y��Xt���M�Ew��w������^1����?����ai��'el��=J�`ǋ�9&�=0���$=(�v{�Ņ`����~��B;g�yR����q
xyk\�-��A,(�[��b]y�%�xF���))��6F֪�es��A�pY:Ttk���(	�8ި) kc��L#&�bû��3�M�;�\��P�l~Dǫ���-+w7ٶ�$�7QX�ɋ�^��_�M����./q�LD�=AЕ\g�8`U�t{%\7PO*�w�B*��I,0��S�o��V���p�,80[���8> ��\Q�묉�U>UR�w�H��������9L�3��F�`-���;E�d���q�0���jƅ�K�d<4��^,��Q1����_>t��Z�hs_��ww����=/�s<�s�B^KP��И	�q������ wb5�$b��0ˢ�ǩ11��\�(�����;�;]�{ʑ�5���H<8�T����]����]�ч��oc���_;I}�e ��Pr�O+���R�|�M���g�+��m�?y%�r�/���������� 6��������%��{Đ"��a�_�;J�On�x�����b��?B�W*;���
ñx�5��d�N���o&鑟�h! ���Y��UVuY?3�6��&�
�\/�Y��o�g�Y2� �� 7DJ�γ��r
K��M�6K�|����F��ms�,i3e�T�j�p �m&绩�8͵ fe�eq��W�5�e=�<HX���X6Y� N�����X�󼧱ay���uH����-�i���e����q ��g?�w8����sI8&}���~+K�m��0M����	��>��\��Td:�D�rw�{�N��|C�����hw�����Q��8��¿�A����Bq5x�R8���N�l�F�x��	&�x�z�����_z5ʉ	g���:n�j}��$:*9
�,��
qp0���K?M"�g;(e(V�:2��]���-wˡ�����j(�e ��dw7���yR=Q��2���t��tAx�5Ǵ���ht{��(�գ]ź�}"�|3{Q�.񂤜�{i��%{���{Q�\07��ۨ=˘$ɵ�<8��P֞e䊼J�����G����~Qxׄ���o]!gq"UV��1�J
\��*���J�C�����0��tM�+��dw��X�,�����1BC�*F_Y=���D�p�-Ey��s_�nI/�T�~B�L(�d��L�(i�Dor�HY^�=R��~�[�v�)_{�}0�X�4=<���[�K����������v�IL`��=���i=W�.#��V�� ����K3x��r�{��tew��Or�r��~&e�'5�|8��Ʊ�#�b�3��=nz�j}:"aԘ�[>
zqt�#{(�&c�����0�K�]�&�ӋN���>:�#�.043�F��ט�J��]�I���L�Y&>9�9��^���޶���#� `��a_j��o3����T��?F�3�LAAqJ2kr.�t��7����W���R^m`~
Lϔg��w� K���=<�3[�*�}pn�p^�k�
��Q��;��,�Wdv:W:{��]eR/s��`���g/qs�P�v��Cfr��+e��9��͕y�=ij�%>��
�l���d�����-e3��/����2Ve��D�
�5{�9%( [Y���S�&�?�U��iʼ#�xBV�߄L���\�+iD�DlU�Q���,���zE�����9RLn.�_Ӹ�HP�?V�-��UK'r��D�X�x\�B��J�GpISE�>�Q}s|Go=!dH68,l�c�����=%;��ܳ���Fr=�	�����hr�O/.������cc�{H�&�	Z�">P�y��߻n��;��n��>�=�=���^hJLѦ�j}α*��x1QC����ܙ��P0;:`�w������Ʒ�*c7>x���ᗭh������ؾ��H�H�3qt���Sܷ2d��m�9�R�	�D��=�$�;L5����yuIQ�e�*�����YaY`q�������(��I���-�'�ido�� �1�O�A�r^���b��6�C��A�k�Z~͘m`����Q��ƞL��O�C-I����A����n{.w��py���
���f?154�j*Hr���(%͔��^D����-ň��Pm��1ݛ�����bFŵ���\{y���1�T������/8(Ҝ@<д0LV}}�EmZ��U�쾆��Ϩ5'd��ѯ�r1�B�F�rM�j.���\��]�#��y�rL�6�|��(!<�s���/rtr��F
Bdc��}Rfph�E(��3��!
4��o��H�Z
Ď��zM���g�kä��d��v���Ѧ���Րoݏ���,O#3f�d�W�X��\�/!_� �Y�hE����\�XCj�NꞍ��k �8� ;u�t��G9;�b��z]�g�I�Rvf����hE��z�n�o!��W�]����R�Γ5��9zF֐��G��2�c)�0�`�h!�*L�X}����gg��_Ó���Iy��$Cq���mB#e��U������e2�+Ӿ��kN��r�J�ә6��ۭ�)�x�</U��$zQyA���)�
|��-���/�z�rb����B.M��ȗ��s��$#3S\��T)��ehJ�����7Ϧ��p{�1�-R���|�{^�G�t���N�~Q�j>�0qy�+��'�Т���
(]`���o.��*x[$<M��}�L��HF��� �MՈ�*�6z�Y��6����W��8`Jm��tp��R4��T|��QP�6����b	L���/�6�S�+!6�^\�\��:-��S���Mlf�k39����Kv�IH��ys����4�͢dc%)B��?�W:d�\�ɵ����G]�EW4�݌�{'8@F�R�M��w̾�{O��Nɋ=B�;]��,�1!�t,i�{�E)H�ZjH�%Hг�MP(������6g��K�ܙ%q��/i�^ܤ?O�;>�H�]&�W�����Vʔ�4]�;� ������/�V����h<xX�f1]N��v��ϩ�^ٰ?)���y�v�����Si�AL��k���Au���y����@��GU����@]�F���[x�rb��Pn�hȬ�46�f=�"BWLgV	�!��X�N��8n�,�ۈK����G�znQ0Vw>]z5F�r�ӃY5:=�����ʙ(?:3=��ጺ-���u3=�����_�?IJ��8���&t�E<�oX���
GO�ürjE��X�=��j�	T�c������WAz�J
�;�`��25���t��7��b�N��'�3���݄r�u���Z}��Q�2#��]if1!͆�so$���8r�$γ��j/�8�1>�<��]���вkC�k���!�)}���0CN���l:܉Bn�����H�&n���Ҋ��p'm��bS�HR\����å�~>�Cw�^Q������L�b1�P���:;�d#��W��:���E\h�:��[�U^}��E�B������S��,D�0�c������0v�/����м����{(3�����!��3#�ϯ%�	%��
pHsQj~�@��
�B��M$NT4��Q�L����irSXN�s�v�8�ʻ*��?e�}�x��Ŋ���7�!knp����kxl�?�+�!��ط���dfT5̎S��^"��8�`��< �K�0c�]ʄ�q�V�Y��|��q�;��x�~[l�
M����O�(��&���'׳�����/�λ����ج�L���:���)�!�)Li�}�b�ħg2[vZ�&�Lو/����S䢖��3�Jc;���'�۵�j/�u�m:m�yzO�~��~$��z3�<�Rɍ�5������GF�?K?Q �Ȣ���n�������u�vM���*f8&�����A�	
�4�j��ڿ,��(�3!�`(۳��/
��C�Q{�!��f$�e<:���)�[�>��f��>Iw�;E%o�)$r�h�	����$��榛�:���lÃ����T[�;+�]T*�˵�F:�E����?g`5t�����Z�ɴ0��+���u�8]�� ��փ�=��ew��<�V������D�!�BPl�g�_��T� ��A�BAaƥ'��*��f΢����oǧT�.�����g<���l
�`{�@�-֏���&e2�a��lGn��x>#����-ݺ�7}�G�w"�j�\��vP��D%'�Qz)� J�}9zZľ{3�1�	�6�W��C�����;=.�>�ϩ�������8GO�m���+D�6t1Z.��:��4�j��Xr㕛6N�MQ>7>��B�$%�)f�{�)��r�ٹe��[y�,�����L�U�OF*��Vie͔6��C�I�;��ǅ;��:X�W?l��ժM���e8�U�kN�:I�8�)1�Cm��^��}S���S��ȵ�]evj��z�ߎu�rƒ��-�
�u(S4+L/4�X@����ꐮmb".>� ,���i����g��6u�fvh���m�0�z'{�cr,ӕ$Z�cM6=������*&����x����>.XY1B���R2do�}��R�rx��g�ݫ�����m��y"��{�[a�*�8��
�:��q�X?
���ƈi۸���E�ۺ�+@�����>��<8k��&��vʆ�y6�����SH���A����������S�a�h �	���,�SVw��'F�k��罄�z3�	'�O�� �"Gh�o|f�Z����m=�>�(�WM������rr�_13X�|�����"h]ָ���owM�dh�pT5�p��隦�����q�<�XF�BԢ���5Jd��z|p�4OH�x�Q�Wqy��S>�����h�x=�zi��˅�h���������bD�DP�L)@=?����(e:���"j�*"�,Z�e�<of�5F>bi��FOਈ�t�!�3��M{zJ�\�`�:��w8��fd �,;T�&K�P3ER���8uQ��	K�F��,�&:*J~4wd\��PCG��t�o��P�(z��8F���K\1�P���(3�2��BbW,��B�M�D��������P���`.'Y��Ɣ
W�e����3y��X�x�c^�M�P͊���I���^��@�St8���1�x�c�L��B���u^ᨰ�l~�+�Y��Ӵ21�b�C3�4��'r��:�'-�ǥ���y[��on�Gƫj�����z��o�/�4	��mj�*�0�8;SC�������[�uk]�˻��zKaQ�j��dJ��R�N�S�3�a�Q�Cmf��Yc<�ϒ��i�g���i�V��<F��^n�%f����ߪ�@=���$�4�U|��=��Œ�mT�b�������ܼ97����hc�v�B���t�����GTH��|dZ����	�8�I�&.+�����>�DG3�v�%���ީ��b��{�����T%;p{�C𮯦/����Ҹ����<�l-P���L��N�����5͏e���R����{�(X��`���  ������o���c#����3f C�B�K��k�F^	z�N����[L�,�-*�
���|&�f�ޞ�'��pvR�~�WAE�F�VV@x&?�/4g#�Y|���i#Z��w�?��hp9�T�R�Z E8������AW`;��[?&�"%��@#C��0��΋�1�{����n���&���t���B�ʍ"��K�[U�)>?�k&*��K�������0����S�X���[�=H7�����(./��-�#�	����Se0�]|T�xnG\v��l����uV"d���@�5WP���wG �n��2�k�Z5��r\��x�2p��P[ ��������\�'[��T�ꚁl����H,7_r5���m[r�>]
�H�U�Nh����0�"M]b6�/�Iء;�����==K��X�"BK��<\G'��aAz�0O)-��1Z�7�\co�6=�bi�=���	��RI����G������y`~�E#ng����5�#m|���$�ۏ��!���Y�X������fp?X5�ʊ���갰*i�]g�.%i�_�Mֳ�|别h����/�ye<IT���l�}��3g�u�����GЊf�����%_u��~p?؆�8sbR'n����~�Ҩ5"��^�̡��O�e�s4��b-&�+I�����]�_�o�щyd/iu;��ۣMPx�������<٧W����tۥ�c�O?'�oz3w��|�X��)Zt���cSMV���lAD��	;VF��p�f�9iSp[�
�BT��J�J,��Y�G�>�x�C��մ~�	:��x��q��
���1RN+j��i��]UJ8��"�'�pC����!�ќ�{suc� }�tm�2��p��j�� ?x{׀'�o�S|�k�l<��'FΆb�*Gb^XȆ���jC�~�x{A5�ҵ��,�9m�@b!��М��H퇂z��*��Ⱦk@�j3h�)cV��"]1x�6Z5^�[P����kV�ʄ�BB��Z����{�K����#׿C/ٟ�I�W�%=:tBo+%����K��|&x��NRXF�y�诵��x�8z��4H0��҅� r#J:�)˷?)H`�#T"���l�>�)�l��U�.@��l���<�`�#�䌀~o��/�����a�5@�t	3����� ��g/O�,�h烈����K�B4�eIQ57���1��(��Y�m�&E�KϺz�R��p�@��� �7W���'ڰn�w�nX�c`�L�/a���n�I���[�(�,�#�bv��\���V1wKk*��|��}TU[j ��ž��]���|�Ђ��	�CL!��Y(Ԧ�wI�Q����^L�o,.���#��x�R�Ɂ��W\�E�4*�"�Xc<�y7Q�rc�eZ��]�N�H�@���v�Xie�>�>k���q�1⠡b����	�W^�R�qx��ˊ���=��e��os�(��6M37:_�q|7m�N���&r�mj������H���N3���%��^4w�B4�	g,��錜��th�/N�^mK��Ar�"6�h4�G��V\+߹��`������'T�ٟ�I��;cWj��}�ve�=n.E<�R&�^&q� ;6���gO���Ię=$H)*�&���a�ȩK$mW`Ձ���޸-����u� ;'Oowyllٱ)�+���p�Y�j9Rw��Q���Icu3>Ta�K�˰���v���I��I��o����
���h�Ä�S�o�>}�:�^/�c�b5��}F�?����Ѷ7U�����E`�:���j�>9M[��ȒWoFC�H���͉�? *b�r���⇖'��v*U�L�)g��[��o�=����z�~U�>6�G�̿���	�=���LOA�M��k&��r��e3�s�Y�<�}��?jT�7�l�dpÂ�<��d�c�?��v]�0��qӖ��&��R ��j���4�ຏyLư���$�µ��63����Sm5����R!���t�ȃXt2�=.s*�S��G%d��,5?�S/�72V��R��_� n^��|8.\U���#�{{j��"��S�P E@�o�P�:�3�nI�D�XD�9#�/&Ў�_���9��PKLZ��?��Ed�fO���l@Xh{��d�o/�B[xZM���2e�1w66��9&���L-���B/s�bF�CR�T�K�2�K�	�v�dmf�[P2���.�7�Y��
O�#��x��)lc/+�}�A�O9��f�����$c��b�g�y�u@>�cJ��Y�$�ꈺ�"]�z�N��H��E��S.��p]v:z�n
�&4�Q����_u�=>@[�y4~��\(Cs��t"!W%P*QPXTi�Q)��� �֮�q<;Os�_�~��e����^�&�1 �9r�g?��D�����zro���k��$Y���z�+hH;$��b�mQ�ޟ��+�����!n�oJa��"r{%��[Z��-�G��@!LLH߼�AV�Q��Z��ع��f����s�.�]��䏠�L�#%iH Ж�	[
��S��Α�u6�=sVQ�ڰ�qH����ʚ̿��l� Selo�-^�b�����L:Q��l�<��,5��y��Ŋ�	'q�v�c���pάj+M��>�#�^x��z��֖Pb����PAQs���Q��wǲ:�jQ�ov��_�����
߭hq��@��CLJ�t����TV_���<��/���5���,1�ӳ�W�]���,nǊ댭��'�f@ЇE������ΘеI���XR�p͖��,����;����g[w#2�۶��n������؆ �!�U�P?U"�]�xjodecK�R����"� ��tx�
{j/K=�}�q��䛝P!�hG���."/O���Q���Y�]l)�w��	e��l��`�UՊS������"�y
�ȅ[xg����V=����L�y`A�#C�v�a�8���_KX���m�z�ӴMت�P6M3�f����o��|p���ݳ˯��%�4���>�>/���E��=�H~?�8��Or���_�����ض��٘m۶m��8il۶m��=�}����?'����<�̼�����1K"=��B�4�;����ƛլj���tK��xP���+:e�(k���q�ws�U~N��?`rf�y��Rʋ[�%c8���G����\�aۼ!۝R����>WV*F��{g�V S�<�,����&iܷ}B`�	j���!}X�k��^�<����x�sr��s�A^�}G5U'���Cne������cE��==2���e���7��s�X0Tt���G�_�WO��'�Sn/q=ۦ��ԩ�]��5��=,p2Ud������?�qHC�:�<:)����	`��id�Ibj�O��N��C��S���������[��x�zT/%e9%�� dS}#�#��ΰ�X�;�Y�\����5����Na{j�5<M.D�,��6�x����ݷex�^@� 85Mzד��֖�G�vf��M�-T�3�F�Ш�U�F\+�i3�F��6H@|Z��cV2���	�?:�����H<�t��z��^�.rZ�֊ȶ��&�sшD��qd���BB��3��4N'J����ĵ�d��B�9�P�����9_��+�4���z��v&�vG��$2=og>ٸ]Z�9��� ��W<|�풫(n������ �R�P���l\$n�{��J��#��z�kqa��8~<m����*���C��ٔ��M��rC7����c��;�+-HU@����8���$+��%',����;ߒ�������yUgу���{D߇M���f7�z<ʫ�AZ��qk)O�A3P���	����i�<�9���O�&�9F!�V��@y������V�5�������i��j��ԥ�5 nN�����#jA3s��]Il��k����Mm����ee�QU�~z&,:_��p��;N+�p�
@�RVCg{:sN�k�&�����<��,u7��ZH�#)����|�L�~��~A��.��Ղ�R��b�߱ߺC�+�e__;8��q��� ��}�ވϬ����D�,ꪆ��&?}���< N<)=���隍��3W��;h��C L9,��oe���$�ڀ<�sSV�d�)� ��Q7��|����M���y�_��z7���/xq<ڏN	�)g4��\��^;0}(�}U<�T/8ȄǊ����{�.�$U���?�`���ٵ�ےnS���g�ǿG0qpE�j��guH���@�<t6���/'�:��ΐ��Q2D�7�a���7����^*mpp��sn;������.��d=\�Zdd�}��~w��h��Bu�N	�D/�K!��َ��My0�w`�/ �W�Ӵ<�'��7��ҧ��?�@@�CBz�x�*!L�}���0�r�q3g%�hG�P�Ҫx����uKH)���q�r�_��ܼ�R����^�^d��G�,����M�=�!�n�߇��_D:�ɝ;��C  �ng.oU��	2G��y��$��W���=QfbO,��د��}�U�t�Q��<����ń��	�A*趩���~��=p9Ar��m�Le�����EO�lh��!և0�;y�
Z�ν$S�}V d�ͫ=���r��q 7��U0���`Y\��W�0w�rׁʥ�EZD���-CM���F�J6���A�B�Z���;���
�ax�i���C�]StFJ��mt��c�}!��r+��8D���ω�W���S;�`^?mx���*����M n�3:�ڂ���O�]_�.nw�աY�׮�=�Ùm!1��Է���mQq���І��w�4�.!��agB/�10�d��j{!n[�zV�ZC\��r���8�?�eQ��w��qR����ne���(*(Fk��F1���s��@3!�<>��tܳc�v'�[d����E���١ދcL����s��� ��EqwZiɖ�j��	���eJ���|��Qg�Glm��@ݳ,���W�����D���c��{�q��5?�L�3��W|6A�x�g��?�����<6'����WO�4H�D��0v!�}��s��C?Us�� �y>��5�b@�����DpJ5u��ͯ�6 -���S��N���h~����k��mtQt�AX�@/-u��T�A�mU1���(�{i��6 ҈6kZ�[�SE�Gs#�I������4��/X�r�nrC�����=���{D�.��o7U�[Q�~D���Q;�ȶD=�4�z�d��ܻ@%��o���J��Yv��6��2	�TIE
� ��p)<�&n}t�4�S>�M)�w����½sWƖ���ٮ�к�T���:�_L���F&�/l0�'�rb�TE���2k�<���^���8N�����b�s����g"v4���jb��O�A�so����5[6�7=�ڳA[�͏e�_U#���%�O� 02g�XRZn��;�.�W�ZU��>PYM����ς���� ����N�S�5��T����lP�Q�x�K�)b[M&^�M��F�����e�P"u����>� D��u�"���}wr�������KE���Q��PR�~U���k, ����!hX8X%+�a�Z�`�f6�}�6��q��V��Sf���}<�i'�ô(qе��-��O�
���teKZ����]�`(y�q=4�+���,�Ɂ���F�.�����d��f�e�}[�'儓M�����N����_����A<_m�ܝ$��ʚ��㏁G-�� ��$М~��@��4�欛RR0�G��K��[�D!�־F�@�Y�6�S�J6�:�&�L��Zj�Nz� ���@���n>:tyHa�ґu����r�gZ���󝮨
8�%�ț��� Rc�����mFQj�עșQ�Uo����j�>��,�z��}e��8�xL""��k��G��F���v�J�E�VH�;�%0�svr���7�wF)���e-~��V\q����?G,̮	�w�J������~.���6���[�.PW7����bC�3�sPCr(�
M���՞�*�t45X81�9Uu������4M}��ނ�H�ŵpt���oV=Ww���tc߉�Θ-�d��^��T��a.��G^�r���h�&�|����{��B(4�T\I;!P���H�A����[Z�QJ��*��I�#�+@_���j6�,��H2tE]V#�Amf�+!e>�-'ûv���8��j�G�qM�P͜��=v�R;k�P�:i_���IvO�#M*,mpᢞ����=��J1��6/�K���y��L �jZw����w����$�O�N�1�P�,6�@�v��p���>ޔW-�jCB���;؍�{*��kP��EW��]�Ӷ�%�y\�WSQ����J��R�(k`�p�7����
�`7)>�|'k��wy���Zg���N)�W�"��~y�����r/�ӱ
s!U�e��~%�jn�FO��t��hL`}ܚ�t=���$=�ɛ�����ɪ{��Y[���K����U�Xq�V�q�>�g���f�O�t��1��7�pG�;ik�_�2�A�$�?��rײ{7��¾�F"��i����������;)_�Zjەݛ����T
��mG� Y��GU��n��s�d��n&g=�/� E��H�/���Q9K�O2y��c��"�G@\M�3��YGfאUK[)^��F���D�aZ�.�5tC,S0�g|���3�����V��FI��0�3{~W�m$r@�����{�pG���!V7��џ��ʹ�̾�H('��^M5�;�ь!�V]~k�U
�Ѽ��
�{����D����Y��Qy�w��s��^^�j������@����g�c$�~��Q��6ot<��B5/�x�NF���N�p�ͥ�kw{A��"2{Ki=q��p��'V�]�$���ʈxzR��v������{����^P���c�w�X)V��-���Y�z�� �G���N�U�Fޅ뗆F��̥k�TV����M�ۊ���DBj��{6j��Hu�u��꣦"2�M6f�ݵ�O��W@q/�DN�Th��=ޝ=ό!�)�	"2P����Iy[w�*��6��2��Kz�-y~��Wy�MS�VB%cъ�f�<�$Xd�H�~��;���n8Km$����+F�5�?M���$���yn��xu哲V���[�����v���5�z�<늡iݰ��Bv���Ъ(d�~k����܋	��]��tS��bt�k�@�zz/6��B<�{0n)����F�5��j�� ��{��f����6���|�����mՃ���F��sFr�2���&H�c��u��1����c'�ď�hC���smU$'���
�{i[��͕	��޹w��^���3�#�ɫŕ���,b%�X�t�Xk�6��|w_^���h�#A��H��{��!��Fc������6�u��ҵ�Ib[�㴔T��՜2p� �ܳ���>�v9��pYKq���)�.&�ֿS�{�a\ExX�Q���k��.B�p54˹�Q�`M�A�EYP@WB��.���ܘ���MuksIÂ���6&�������)���V9�i������j+L�5u��U�B����}W�j:�F'&�g�����ş�a7����(���Ƒ�Y�8��#��O�X��,��Hx���e*d ˅B�G�)�m�Ws�� 'T�Bx^��QɎh9�`r��Y���X�`���c����ң�A��)�'����F�ten�pLÃB(I�A��s�aB��=��h�j���#=�O��k᫛E�盃r[��y�$���H�ek�B�\oי��QV1�Yg]�Q'�?�Z!˓,E�����,���]Ӆ)��h�o��RS���?3��Y��mF���j�u���	&����y1�̶��V�ʛl?ܫֿ�l�e-���mer8w#j�*��]m�	"î�&�t��DlS4}^sx5��=�І̘�y��dr��D2�����.�WA��_!!1V�0�N�3`��Ƕ������)�K��^2B�1Lgڂ�b�$��s��|T}��m��g�z�h��� �^i[B��m��q��I�t.�m��8`4�Ah��p��� �x��n.�w̃��?&9��7����Z�k��vх�۽�Q���|�SXx �]\"���(����5��?EW�ҥ��o�벖P L�`�����P�rL�7��)�B#
ɜ8���
�o?��2��7/�j&�%����Je1���P��C����m.��?����t0A~8�!uƵ�A��A�1���]�S�_L��E��L"����:caay�\>�澫5BCS]X������P!i����Oj�<%�6V��j!����zx���0T�+���q��|`��������~b ��E	R��:�/~�
�i(�xGc�e����<o�z͢1�$޿�{U7��yU�Mx7�n�5��|�"��B�G�s�a������;�vuT\�2�v�)��)��0��ڕ<�W'�2��2����-�C_*��b���p\mt6�������B�����qϰy>��_mj�^ �+����A5R��I�h"�Mrv�k;�P�!`DE���ר�}��`0�6<��n?�$�$$��^���2�w�3_�-Z&"�P��3�L�:V%t�� ��,ĳ)��b��kO��;��ӉoJ����[�8��,y�EuF+��#����
�nmAL����g�}�h��[�^\��
_˴E����Q�����+���'�h2+k�eZk�����;F^��k�{z��{���@���&K�hϥ�`ӡK�a����K@ߟ���ZՕVÚ���e;��yK�=�h3꺸�u��3�_�S�Q�B��k�LT�p3; T���g�#�����L��kP���/еj�m�����o6�0M{�I�J$����![Lh�<y6�	��D�e��#�v?b�'�R!x�x��=v�休���uL��X�1�b�u��h�2Z�.�\u�nL%��,�ʦ��·��#y��������/��HH�Uy�d+��V��h*p���iv8�C�cxyI� INI�H0԰W�g��$p7����^�W�����l �U�=�q�Ʋ�Lu����KZ�{JJ���d#�޼�j�^�2T�A�:Z#AVK Q���C>Ϯk�K��] %����G�{H���
~wݥL���k��ۈi#E��<R0���mByKO��D�I��O�jw���!��;�Ҧă���َ<s�Aʣ=B�/�|'�b�Vh5���5�ͤ������]?�k�y�B��C_�q5Ϣ�g�E/n��F\�<>?���8�ϙ�z�5�9�����5y��1Y���[��o��ix|Z!�N�'�tn��%:XesHc,(������Նnಎ6L6�(�)�~�(��9{����G��]j9�B�z�[�5Y��{:I���׼qHL��UU�A>�>C̍
�T�k:���J��*\)s[��fl'Wh_b~s�>���!}ܺ���������O���l��u#޾�\VJ��hK��Ӫ�<1�j6={~u�/&a�;&F+}/��C��O<��0�����\rb�di��I��3�Ew��h���{�יY� 6�O[�lI9��QQwҌ-��ːd~�{'R�-�_�x�����m-D�D%=�B�XmKv5�O�⪣�FB���Q��jE6#^ud���9q����c������7��y��U^��V�]�����O_����Y�?ˢ	�1:T��P(r>�J�w*�H-�`A}�O���Bf+�$;L''p~�Hj�sm�7`'��[|T���-F��$+sɗL�ʣ�-R���&j����Ik#k�%Z\�+B���^O�Z�<�t϶-B�1�3!Mj��]�K٘������j���txsB
��r�S)�H�s&�t��O*.�A��Kb>d���S�M�I�\�����n�G�q���u0��ЊfK�����$���H�����4>����)ڟipBV7!Ѳne"!i��xap�:	+h%I�I=��O׈>�?�Z��~<l��^"(ε�l�ᝍ�*����JN�=Z33-t0ã��Ye�Rփ�fn´_w�c���7q��lE�G|Y*���	�:�Zk����]�����Ji�w��ǌ����6?�?L8y���ݵ���'jO���=���6�x/�i�ڛ~)�G�VK�BBҙ?��̀�˪�����E�.���\wF��	�1j����y���{&DCLDQ�������x[�~�pV����x���5w���K��pkZ7��hϝ��+���<=��sTI��i��B�V�ɆB����o�oՂo��^���/���ڸ����!��������v㌫z�R���?㳰mm�Meu��$Z�7�'{�/�jW1"��~��O�+ ��b�6.��j�~�	E=��|u�Y|Q�`r�д��0N�3�T���V��������V��ަ��d����:� ,��͵��A��Z�׋�i{X5-��g$W ܎�1k"ܼ�C�$
�Z
7R�
=�V�ПH�:�����r���l�9>�����h����YoR�@�l+�SlD��{�zik)y��@>/�r���-mu_����N��lgc|���K1�6��-~�D �EOG]��~r��\!jd�.l����sc{P��9X�3�/�c�	]{Gc����*���L�Ŧ���?ҝn�\�>MxۨyO :�-�ۙ�04������:���o�D��m.Dc��&�m���!��������F���g��4��\���ls����6h�L�]��"�I���@[���n�:'��n��}�d�\H��6��Xg�c�m=��Y4G퍶F����ȕ̠Ҵ�̷��}s�Q��z��y]���Q�V��:��E�t��"�56��-> ��f+��q��}[bd��s�t��zl|�7�٨���e����N�[��^Sq�$2$��(�v�]t�/�!�_�A
$a��f�c������.]��:dσ���T�����3�+�Sޟ��b�۞#��8�Ƕ'`G}dY�w��Cw��4��}�Qa�z�Y�צu�����<0�z��C�m�O�Z�uQ�u�@��9c�8���ℹ���^�^�&��*Nw�f���6��p���O<��.t�\�ޥ�b���IkG=�[�4,J��ͥ�B;�j���d���+��F�o+A�X����Y���Z���RH��`���Q��K�dG%~"�Zբ�V�9H��	*���q4�_��YA�pC�]��_\�$Ǵ���f���n�a���0S�T3f�Zᄾ���y��̊�pպ�!�O�eB�4���慀 �*�w�/o��pG;�*I��d3�k��]]��Z7jk��|'�����F_ߚJ.m>C4�N"���w��!J���&	�K��q�����-��혧����ǫY"G�]����d�-L�;;&fyru"<W")`cs������y����d�vs�3���GthM��ի~4��Q��1��e`��-�Tg5b�M}������񻘍τ�v�P=j������V�D|�NV�<��N�[[+�����i����nk�X��[�N��\��c� ��M�q��a��hÿ�"����d\>ml���|�>�!_i���O��F�⁲��Ы�j
�� ~ً����>0�1��'������hY��|�r�8<��˛�R[y	�q6���x)�_eUHjU���I=t���|^��e}2*��_���$ED�z�}b3X�@kq[�{<\�H���ƶ�����1T�
�30/��	]Ԫ�:�,k�~���j����n�[ݒ~��,���`�e������Jh�\�#��7ͦN���ޅ=y���/��?���o+�+�?���5�I��ü�p�ԙ�/�|*c�)f��HK/o�74��@Yr*Fr��e\��m�n�]�l��մ���Z��f��7��>j�j3s�dO�De�c�$MS�:�,���ͨ���&Wnd��n�L����� w5�w���ٍ����M�"ȍ�^�ӿ� g[�w�D��׋��ٶM��$*�	�2JyY8+�
[��o�?7��	���ࣲ+��@d��@�U�i�E�9����`���Oخ���ݑ��]��˥�#��0(��I�+��?�-,��jX�1�N^U������'k������D��3��ǐ�l��~�k�]�d<7��)� $yʓ�et7i����6��}Q.�r�+sҌt���<Y8y�zKObw���/׹��H��m5Z�χ��yrp��1�AzT6��$��w9������z|^0xGX��˺�w���멢��2G��֑�I���dn#"�VO�o\Hw����I�ހ���DZ�@%L��'�����u�����&� h���o&CF)�}�qd��TŰ�z��_�p��z�_�僜*��r��'����m�ϰ(����K�o�������2����W$�'�3�LB7lğ�BMf�Vy���rD
��d������ޡ��R�U^~��QX�\� `��pp��`O�b�t���j�E��¸�1�?}]�~���j��6T4�5�(@������k�o�IC�Q���Szg��H,��,4��ү�<���!�$l 	$#�ʰ��I1ߞ	@Fwd*�@\=N!���9��� �i��a,����J�J��ߝ[��@7��*��6.D�F��Y"��P�E�ܐd�M�7�L#��<[��3e�N"��u7�ګϪE�J��+ ��M��e���V�q̇�6u��8�9��R����<�V��e�{�2��=K��5�r�z������e����iX��(��Ou�;4֚��մ��M��<*��*f�4�Ziw2�����ĺ��+��4�2�(�ͫ�+@��XjL�|��<������Ȓ;8d_�%�q!�l)	/��9O.��(��W�ǗP�|�y����Ֆ�u@	�!��w�'*���[���vR�([J���)TM�Hϋ�e�g���c�I��b[��k�i���!sl�ᔽ>*�l=���"H���$�W��d���d���
����e$ͳ�\�c\A4��ɚn9$�k׽pLu�6����ƞW�>���QN�����r�)ȉ^r��E,�Ul<�>F��V�j�t}�6��<�"+_W&V�����J7���@N��=���A���t�_���02.���G��!�nɐ�|:O����T8�(�+�E�)�z��`�n\&��d4B�G��w��~��T�����=??�d�ZG-
�6d�zO�/��~���B���^�n"6N'���������X~��֟��$�z�6c��A#�`�Ɗ�/�2��4���m�Gc�"%�@�|�]I[�6TML��E��7�Ɲ7s�������|C�?=^5�Z7ļZ)Q䭻KQrP7�1n�&�z��?#�j�q�4���U.��O�zt0�g����S5qN^�O����k����m�0�;hR����4��h�i���f铑lm��?/�)(��2�oE��Я�f6zy���eH��e���~`Rr�l ()�������@L]U	��MƕLN���gbNE|����?�$=h$L���0�ej���;]���Ŵ�v�c�<a;�u;�1ˁ['�y3_���;r�$�s�]3p["T^��6h�X���������x:T��)�6^RBI�h���?�,Xb�n,!����vQU�uF/�[M�c��L�U�F)!����{�y��6��D9������LMAĂI��vǶ[����D��2�6ʰH C�ט���O�N;|�X�>��(���7�v)	�_O��`=���!fUL��l�X%I�)����EyO ��������]t�6����Y�!�����/�戁�]t�3�m�R��j�D�T6nz������F/"z��wQ�5*�e[�^�HA7yy�mt6��._����|��3«ɞfcX�C�	����e�B_��&�``��l:BWw���\�[�R������v�_ у$p#�WK��Ov*~��2��]�m�\o'�ymE��W.�ϛF��Eұ訃]]t�͉����Z/D%&��ԕl�g�0eB�nW3F���*{��f���E&T$�q�!p���{�f_k\�/w"V(۔�+&��
�����K����z0�*��N�!���y�+�ڒ����{��:����n����0F���B�䠫\�Z�"Ts�[2�H�O;"�D%N��1D+�X.��=���?���Ԑ��p��1S�L�vA�^Ԋ�9~1�m���j����e�| dt�G���P	%�zh��9�(�(A�=���El�L޷��gsٽ��X�� ���.��F�
<�p�Q]�ˆϏ����̒_ݽC��
%��_�ID�D�F��Y�	5ãRp�3��������E��+�g"��l�w�fvӈ�����	%^�� d$�7��-�٬˩���R�;����=���-��R�E������"��F,�%�����zwȅ���6iu&x��yt��
���VT|뒕�/ yګ�
�7�*l���6r�4�����5�l*�T*H��d�|���$��ME��<n~����E,�s���B1�u�pݵ/)��N���
��ę��3=��O[�	6�j�|�gҿB?��F
��I}:�K*��2>�^%^J���t���mEY c�������S�}-GEF��jqj`�̧h��$}�ҿ��BF)��Y�^�� _�e~Ϝ`�����ѓ$�dJ��_z؄���3UCt[����o�F��ض6��6}���� ��s{ =B=�ߛ�����ջ�-K=o�H���#p����<�*W����$�H�^�7#���E`	^��T�^YxT-$)�^��.�Z�f�Rf�F,/t/*8o,J�H�0��]<�lig���g���#p͙E�dr��bz7#'��WV�OZ<���<2l�K l3��a ea}qu���}��d�]�y	 �_����*�a�#KE&��됣��z���^[��&&��<�1��x����A���s�"-���O�:<�4��f�J2���l���>� Uqᩌ|,��c�t-@N�X��������H�^��b(�_�����B>p��l94L6�>J�}r��8���k�\㉕�@�빚�ㄏt�`�,B�3A7�U(5K$4bsOX<�aI�{��]5E��8W)*�,��}I�%�t�( �}�_z6���kө��L���c����O���%C�T��?qϫ�w&��I�:S!q�\������~���Pi�7��\X�ns�S��Z=�$�y��<.���gs�p�k�F�_ G�g~��n�!Շ����tgc.'{�z���>`�<�X+�0 �8-
\� �p:/zn:k�?t����E�!#���iHS�k���Ϡ��a���#�0Q����A!n $ǡ??��`�)ުX��l�z���	��A���n���=`��N܂��-l�ʩUzr֠W�����������O���S�]Z��!��;��	y�۾>I��cPp�Q�֐K�f���܍nzm�qk#,�ֶ��Q�'�ݓ�%c�������H�+%R�Zo俞�.�r���n����*̞g�[X��V�)��a���p�i�A�:�U�%�zSm,�3�]QM�<�끵}J�DLM~*h�(�rn k�K�i��Θ��	�f����s�sCg���
���Y>��^�g?���� \'��ĸ!������j)yQ���J�~���<:���It�ܭAm��Zz*Ù� lB[͓
��_��[:�tO�ǜ}��_�^�8����%F����{��z���[y�*���TKY}�WF@�*�H�?�T�{�y��M��t��<����o}��"��λ9�sm|�1E���'�E��<V폠{$�v$檶������.��x|u�$~)�>+��=M	+VL�J�*��f�K����%������ve\}1N鄮����f�r�D<�ag�ZO�?=���Iv�c{6��V\G��|k,[��w�.�l��Nd.�
��m(�#EN�b+�K=-32aa�(o���2�KJ������u�H��k�¹��B��ܳ�j���f��z����°��F��w˵++�U�!�(e�n�X������q�\<Z\���no��H'"��ܸ���>??���ĵ�C3���4�0�Ͻ�ɀ~�T�.Z�6Y����or��I�kD$s&�@��g�a�j$��+�L��BbqƦ�d�w;p=hӵm%������4�
��h/�B�Zs��V�p�~UR�\�|�����◵a�S7�Z�-����Yl8��bzq݃�?ՙ��ƻ_���K��Xo՝����}$2�ء���X%��B��R�ᬪ��Я�*�w�a��{��A�;]����zK���W|#I�	黳�«v���(y��pڬ��Eyt���3��fmL�3lC�����sޭ>q�FqR��%-a���f܄�"�<-0 W�� �̹����g���� �k�$ޭ°\ˉ���(���ǣ�x4�;���ePgz��,'��y�.zY�Y��"޸�O����Yw�pG�F��>I{z�ZL�����|�)>^f�O�t��c)e�le���C�h'Ur=h�hz�%`�|�<!,�D�"C� �'�7dM�7&MtY��T�I��7�䃶�w�����Sk��J4)���~�vG3e!hu�ܧ�M�����&ב9u%N8|�%RZ{F�"�M��9���m�V�!$}jZx�9�fX��nP�_�U%�h|��5�g8 ����W��յ"k�h���'U�o�+��|<0�V6�ű��
���/��� ��m��P�f�^�����םP���n��RA�pR]���:t��n�������N�s������4����Fq�)�GU�ۉ��� b�/S�RA�Q}<.�f��t���àm�S}���VPr�`��(;]��x�8qz&X}�	j)�%�LVN��א�'u;���;X��7���l��r�������5��c�@!��T��] �%���A�,��2������kK�_�U+�R��}���!C�4A��e�]/V����x��+A=�pwI�k��s��>r���{�Ű���9ө[@OAE���~�˱M^4�$'�|��C���ye��[qi鷒c�R�}�������,�q4�m�^r�1i��6f��^%p���l��!-����w��lHO��?K�C�Z�;Z���A�d��_n#ݬ�[�[&31C+/��+fӮ�,�Vu����k����Z\(���e�3A����������>����\��M:�,�0'���t�(�03?���O �������uuc�^��(p�8�����c�K��\�,{�N��W��� Z��".ȵ0`�^7���ύ�v6��VN�0�x�8�v��]=�����	�H�d00+۟�3?1^gh����	�
��6�]�N��W7k:e`&q���,�)j�d"���a,)�nƩ����1qK�%˻F�6����$�q�"V��ab���\��A�
��*;~1�ܞm�2R�}qP/�Q ��$�'ci�p�4����X�q��G�R�W����\�r�����`�2og��R$tĘ��4�jO���Z�*�����-�A#�ˁ�����/ EW�ه�h�ric������t���ݰq����}Ҵ
���n:�#�1��X�g~��a��Y����P�:'3v
���-���v�������*����ro�""�$��{��ݦQp������yl;911z�NK�MyXBi��3>��n�K�1�g}�UV����m`1����[���s�=X?�+i���:�n3���T�(w�!����Lķ�y��Nݥ"m;\�S���u,{�x�L^���ʖf������j�#n��e�����}�ʧ��u"��'*Z�x�
5Z�N1 �2��*���joM�f�̞
����\�^=i]��.U2��ʲ��{���vχ���ه����C�ُ�z�H��,M\�i�Iw|��"G��TlNR4.���������Of*~Q,�+%��<�����k���b'�����N3曳���"�����%WO	�IVӑf����}�����C_���ï��w�
�P����h�W|��b�	�q��(�g�B^i9�N����~�V���W�_�)L=5^d��+|&@/���>n��Z��\����P�%� �Gn���YN䂱��5�ڀa�d���#����[��M��5Fm[bK]B������\L#4h^��P=?T��*0�yk��;VD��4vE�
dtoFI5��S�5{���{���/$o��̹p��Fuˆ�2c3��n��s�#���\T��6I��e��Х�P�X�6d�ۃ-։[v��S�>Tz�C�Nr�o2.,!�g��i�V�o-�ڛ���x>�>'chV�J��%��f�8膩2
@�bLߜR�����)�d9Q'���ܯJ�K�!,&:�W�X������hΤ����oX��^9b�O���ҟ����*�����c{����gn���־���m���x�}c@�8u���P>܍>s��b#3��|!�r�z2�9T�$%m#��������I�G�����&|���:!P��+Ew"b<X*α3H�9QŸ�����Gv#�&�R��xҚ2�W�e�� �P�>�H1~&��}�5�V9������N�˂�|����Ռb��@�������1S���/�s��"w�N$��T�s�L��2�B�.�9s1v-n"9+��;Eq����&/;9�>���t�oV!>������c��� E*��	#�� £���N��P��:䭺��"�-�0(x6����Fs�,9�vھ��b�C�յ�>�rj�DD�<����YR��'��2`OX��b�&�xy1И#0��Rq�4}����<�4���t4�҆�C���Z\`{  ( @q�{�`�O�(������6V�m�avOq�eÎȋ�NRƲQj�I�x~�w Rԕ$�$�>�dksU��}�6.5��\+�͚��MQ��)Pj�z�̖��ێl�Ui
\�����8O�����}���e�E���h�ach� ��&�?խxˊ�t=�f,��G�ԍ��3���Cӭ,u|J�V�Fc�ݶcE���ʍӶe��D*�u����1$��M�߇�oc|Tp^�.� �`�GY�uǦ�?�r��W��so|��f��~�Fq�.E:%�&P�f��ٿ;͒��q`5l4^�ZR��i���wݡ�H�d�
�d1���Lݪu!�P.`��k(°i<Ȋh	�� �~ҥ���ry��Bu��x�➃g�r�s�Z_�n��21A��y�P Y��y�n������	}/�O~��wH�T��Zm2ӃFcc�Z�4�u�ùf�F��-�R{ͬ�T��E���x�����˄Sc�j����YԔH�=1�հx߅"��lZ�����.�)�!�g�~���ȉ3Q����)E�f���Le�>G\D��ޅ�����j��X˄�O�B'���H�.�n�#��8��t�C�����[GU�v��QQ��m����H�H�tw�M�J����H��" ,J,��\��|�8��3�{�co������sNvߢD�^W��k&5vڎh�ã��=S�+'s+���Gߎ��.�9-���U,	��-V~��W��#&�O��Г}�Y{c�m��]u����Y��Ĭ;�	D��VS���w�F)�j�
�|R�s�7�"����7'G��H�S�����ɼ�q{:�{��@�YvZ�m��+��j�p�t��Bz�����A�ȗ��	�_���S���b��璘��d�_�|$�K�r�~�
�.�7���Ԅ���Pq�A,�x�ZyQ�#�,f�-�in��w�b�ۛ��}8F��6]���v�ٳUS}́gA6{�W6�wV�i��:$��HBI�z�R3��M/#�#HD���o�8�b�s9sׅ����U5�wM�':N��.�r�{���cZ&\���k���3bR��\�²��)Qͼ,�7��HG=����ZW�bk֯�wRcEw�\_��Ř�G����m����ܿ���,�8�kk�sAq	�;�ܼ� {�L)�A�tY͇.K屫4��X��im!}�o����=�[\�(7[#�ϓ���!�#�Z�Q�!����kz����z<Si���꣱m~�6��,�]�=�`GݬQ����U�E��h��O�DȄWk<ֺ�/}&��Ѻu�&ڠ.	p��,�k���A.�X�3��$�n��Z��Ʌ 1'X.���Ď���~��)Ћ�v̼0�,.�DEſ[m*�L����1z�jՎ�J�����!�/��y�X�]-��2>ޒu�CX;B�a��(z��c�"�?���e��~������w+5K��
��ɘ��VL��o�(N�����R~.jK3���H�s��7++L��J� �`S���|�D�iPPkpI(��[Qf)�ҝ4�?�Q���O�UI
� KX.���2$5�� �[�����_��,�D������nֳ��*A�U��D����?={ט��r�zY��ց�����2���uft���������L#�ӎ��.�\rB�qX���g�{}Ò��^�|D�q]�I�a}|�Ʀ�gp�a����lDY(�Gek|�qo�zq��q|�}���?����p?�pj��M��}���>�w�u\��T�I�9��5,�s�]zdh���T�cf�4^�A,����RL�ܡ[w2��T�0�m�̗�mmq%_�d�
^
?��.�''�"�KI��#��1��L�)�nx��u���k��^��1�!���:$̼3'�k"/]l����o��A�7�D�h��������u��g]�T���W����]�[	�0a'tAYEf~ָ���lI�n�:_�m����Y��U�CUG8�0�0!�۰��K�D�~�M:	�E�@�n��G���=7ۄ�鳃��d���<'͔z��.�-՛o�8���͞F ���� I�+z�3��cϝb��(�[���d�e��:[���%6���U12=��|��_Q�=,@�~���&p���u�����s�e�Ҏ�����S���On�V�gbhM7]%x��X{���k��Ͷ��N�g%������l�)w��;�I@�j�̛7�/�`��Mb�~�m'�Z�	"gh��@2b��nDV��178~$�K'�w��d⌯[�/����l:�~��L��|�9=)��/�q:-�k�ZW^�uiZ�����i����X~�QO��~R#��n���f���G2<�8P�,���lo�U������r�&�͊+l(�kE�&g�gy�h��M���\���7O�kA��H�e33G�T�T��.;�����m23�WR�'��%]��8i��DTL"��=OF3~����(�;��\������qO>N�{x}�z�i�sZ˧�.�[�V��^7%0׊2����K��QUvEr�5_�8�'��s�%���w>�-Z�b^�n�י�
o����9��;������8Ǎg�ڳ�]i�Kw�I�+�V��."Y��&VG���Y�כ?��b|3��2�P�娻��B2��`q�@�q�������-���r!�v������8�>i�FQ0EO5�;����M�e��N��� 뉥 ��׶jc�����dm�w��b�Qyx�����rH���B̺٩4��(Z��I�j�ͤc'��闉�[�*�n��.�\��^��bg����"Ҹh��Ƭ��F�6ݥ��_���c{nb��RP&^"�j��0�5�Ԃ���֕��d)��-ն|4�%CB����o���ί̃�|���:�����G�|��������WDTI]IO��U��x95�qz-���wW��2@&l��ԚR����{o恜�Ţؓ�B_�e�q︭d
��O�]��(��]O׫���ʟϞ�_A�+�5�l���(6p�� �໦���e������;��gQx�b��M�n�|a�4���;_���C.߉�=��u�
(����_���)�ul�_�������Gdbŕ�f��]�[������5u�,"��������M��=���?��8f�?�RRI���Qjo
��>ʴg_0�4�/7ո {��-m�G�αw�"v�\��=)��z��,D�dL��8z����WdI�.�MRn'a9���;������^�r�����)�A�1����'V�V��^�Fjy�$;�\mR@7�UcLB!��b���g�2��D�ߟ��x�&?�NMRt���ű"����Җ�Eb�DaLJZ�(# ��IDp;�	����Mu�:�P��ʬ�;���Y��e_������:�R=,Ϯ+\�b�(��h��=)����ƃϡ�e�^��Ƃ��=�F?���W�ܚ��س�3��=���O9�Mzd"-}��FP25.�w�A-��������W^K�Q��lw0q4MO��lwU���KFo*e�jHD��_X�	���^w��g��y~��3��U�$�)�0h*TO��flty[�r��Z��'Ϋ��,.��T�;����W�z�_*���z6VKLr���YJ~eY����*�{�t>�{E�vt}~�B%�����{:r���@�������vJM{&@�Qj�*%fsv�1���Cow��i�*��X��ʂ.ӌ�uS:}B����6l�_���v��ڛc���V��Qa���4�šP�����N�&��5��:��Dky���w�[�z��Y�9K.F۫�p^!�i��[n���٣*M�1/��E��������)_�>~�z2;�ݎ|Я���c�uSۡ��V��7~�\<�Z���v0Q�A�Ȼ�v%�Ƃ�Ίwd�i������>w�R��Xc�c��磷�[	��P]{���IT�TzwVI&����x^M�gߌ�����+�Ի�<����F��$�/|���K�Jn����"�gbК�,��m�Lz�I���X|ۛL���w�#���A,>����h������6U�y�j���1CCeKs�I�)���L�.�����;Z��迷3$����rl�.��يe
�O�^��ϺѰ��*�U��+�LiZ�F�m1���m�'�ЯH��1#`�\a�R߶�T��$�;����MC�u����[^h�k�D�LD�B��E�����ttg�e��u�-D�t��;?��X|3A��ӷn��w_ތl����?�;�^���!F�Ogt�G���f&�6�6�!����7̹�͢S�Gw�;%�����J�$�;M��5s�5��W�âF����y�&��N�G|���� k�K92������F���&ǫ�-Q�v�9}�9�V�¿����V!�vH��Ԯ'z�
�V��g�wG]^��JK~j�9�Y�^�jߒ��v�5�D?��ҿ~{ߴ��5�fk]��l��U���I�����r��U���[���z�7W�w��w�ÐÈ׾�z�{i�vg���\�"o	����V�M)�B�,4�� �MK�Ţ_*-�o�a�J��-�6!`��7�D��|��;�A��sym�4�x�	����'��(���/��(�?F��|{�8�,���u��	9�ӈ�ֈ�_;ːHz]�p&O����|�^O�"��}��-�7�*�F y�ܠ^�������@��6.dCMpx⼝��C7���ҟ/��;~ޚ�"�q�^zi�g��*��R����s�t��N�JԲ_t+�h-;~���Vr��<r�ڛ�tnYv�y�d B��h���v��9�cJ�M@`��RHݑR��%���� 2{4��O���Lz�G�D�����z0L��gco;F�3cu@�ĩ�8|{f�,y�n.�n+��WG;�(��1�p��$����[:?{i�6�o){\��P��:K�׌ƭzǞhw|y���-,�nV���aI�'�� �o�5����l	^Y�g`����$���D�)��^�	e*���4�lnЋI���9q�Gb[~��j����y�J��dab���12�h1�0��	*]<�q%��L�J�e��>z����vz���I����7{�+1�&��]W[��c�R~�&�,��Els�;'AS�4+gѫft�=G���2��1%�J�q�a&p���Ȱ{9�p�Vk��ԹJ#�j.���'B�Q�]������f喢k�z^>d?�&;~�%�8Ϋ(D�
�h�R��}�������j�G�I��g�������<�U���
�;欭�sT��ǧwnf��n{j�Zjs��^hr9����RO�<ݿ��O�(W���~�>��EzQ��ud����+��ܙ9�����|���H��zC���功�iȗ�_1	6~`�A^&VQ��Nc�)b�ύa<���6�>�0B >��V��u�O�3�n0
�]�n�����n�	�O���1���̫'Jy~�e�\4�_��k��v#��}/��S�`���g�w1��v�d���
�k��G�V����2�z�z��lǷ��H��c���% �A�\ί#��_VՐ�%g������-��߱QbOJ禇Hi�����WJ�5�Ó�|��ȓ�I�/�K.g�Tҹ6��u"A�f9����^�4�
��:�޾���Gq�n�Tg7������8`p����ё�+>K��d���.DA9yک��-�{���.�-�0�O����|����V�x-eڠ'f�pI�Ƈ�\����y�B
&�a��K��q�OR�f�j"�ȿ�%JlR�����AFR�c�?�`x�	�4g�Q"uW�|í]|E���������R8�:���8��I��q��+�F)H����Z�%>6�^��!��;�����K�ɨ��&t�.vx�Y��oX��?q\��V���v$��,���(���ذ`�vؗ��ϗބ�����7в�Q.�U��ft�cq9*DD�k3l��F�� �)�9{�e�-m�̇�'�X��@�0Z�ۿGXu��m�׻2Џ��Y0�=G�i�����=�fҢ��f�C�Q�A�.e���̒��K;pma7�f	�5I<k�b�Qx��W-m�������]���`���?�P�z3v��HP����`靲�W`�f�<#�=��yim�XJJ7�gs�� ~v/(�����н����R���U�h���o�B�&�8)��S�4�[�,?��U4ù�='-=�0��5�9���8G�Xx̷�/��s�^��R�*��t�ą�e&i��>������J4�j� G�ҟu
w�]����Z�햛B�z�X:
^J���X�;�,N5bt�*Ƕޫh��nE�K~L6ܿ�:�L/ި�h ��^!g�C|7���ԧ�@��K��M��IFѣI��������)�����_��I�tch�kD�)�κ�����
�����[1ֈ ��ރ���K�V=8- N�(���}��A^�;t�c����!߷9
:ׂ{1o�5�i�m�<��:F:�=k�n^߷�G�>����Umv�9�h��2���X���Zk�[�:��Hj��0���]���L�A�Gg~s2�Z>�ץo�	��i�:��ͺ�ْ�r������3���3y�ӷP��_��V�����U��^�_����G����b�م���n����<�&�Tx���k�3)R����KߑV���㻃y�T�4����8�B"�`���Oo�]($��q��$s>���㛝��3yN�n��'���qħ�.#�������wx��C�T�TT���S�%5��K:G��[߉ ��N� \-�@."i:-�[�k��1(�GG��=���(q���v!!*�����~*�r�Pxmm�k͉b��J�s��
�e+NOx����zo��	
˙�Yk��9�#Q��d?Y�C��бqD2���R���Gx�]���vmQ.Tr�a~�4�
��P�\ّs�fC�ˍ�:�L�a�.ꏄ�Tx�ح���\���7~>f��	�E�9=�u׵���z��3�^��=�F�_��T��	{ ����~�=w�e����/n�'��8�7!���[N�57|txw$S7Tg,��5��s�����_o.�^�*��wh����[iU���$�J�)�9G.�d�y	���%b�G��k��x���ρ��ρ��ρ��ρ�=2� ~2��={���M���(e==F+t^�T[i�/_�G
M�չh�����B���5J�5�u+�l1*/�/]�$�8��"g�ͳ����f;^ٛo��S�����!22�q���h��e����1��ʰ)�����c<#a�Q��Z�|����oߝ�a����#�an�bsr�E�mI�ԉ/�V��	���X	���}����2�pdTT�"F���RAc���J��=/��ɉ)��&<�L;cɹP���c�G��|��r>,���8�,`*���&%��9��L��>�7׭�t�ޙ�*xU�6V�N�z�[tm.��9��װ+�_{-�Y�k.C-�e��nn�H�dU���<�Y���Ç�L����49x��b�k6�Ł��#w�S�C錎����XQ7��Da��p�ƪ��*�t"��Q%{�֟ʩO�]�M��;8f����d��TT�����8l�ʴ�׮G-���X�e<dxN�Ť�X���� 2���ܧ>�b�N�{�wt^�|9c�Y}��-��w#�7W�l�
Y�(Q��_�̖Ka�<9� � v�T��>������G�c2q�J�eZW>�����ݻ�<*]�,����$4Ht�������Z��f����#p��������-����&����yU	ueee�#��6�)���V�w�u��4n�H�[M4m�~L&����+>�b���G�]?E񭁅�2;���tv�����m��+�gS�v��[���W��r�l��r�L:��~} 6����tc���:S$%�x��w.z8ߝ�����e�`S�U�Kj�]:xa�Ȍ�����Ǽ���qC��`*�0"&��`S�pC�r�I�c6e�J�^K�::���;w���x�,L�x�2z��SK�V�H[*p�'�������w�Ȉg�T�[2�Sԝ���TNZZ�aw�_�'Y��@6�T��ňZ7U&����Q�l!�w�x�_�1Q�i�s|�< ������/�g6��C����j�T,f�)x���p�5�u_k��n��wn�"�^�u{ͱ .MB�g^u�:W�$H�g_*�Q��oj�0L��I�e��^bk��<P�y��+G�[�z5���Z�޻f����	m�`���BQ��\(fU��ϯ�0���\qY|ُ`mjjrX.A?��^�{��=���� �^:A����#��&M�$
�dS�d1a|�|��Du�P_�E����Q��-�J͎ڵ�~��`�ڻ��u���LOOSٿJt��v��N ����E����W�N��)9�?���yc鸝~ۘvp�V6�����W��P�`���ڶ���M=��E C��R�t���a�;��F�! 
�)7̓s�7W&OTƮF���n>��p-� ��SZ����O��P�P�7ד:_1���b��l{<#)�5�Z	yf�~�������`� �PF����#�0�şԼ��K�c��"2RRH���nѕ����-n:��hT ��'����e#kE�`�
j����&��!���!�O�L���%O<0 &��Oʿ�C?�AT �Z?�N [5[��K�Q�8%�y������Ge�v�@"؋�� �Do� V�7��e�ܓ���޲�����O���ڄ�Í�p�6�c���ndQ�,�^�#$�qou��͟��4H��t�OA�Wh�,èٟj��m�6�م v��*�m:��;�d/�$0BI�#aώ���E�C�s��9l�������m�W,q��;%���j��3Pv4^'*5u i)=Y�S��R�#'��w�C����&���Ce� �7�V�s3��ʳ�����z8P��gb"�S'77�I}��s�t�aly�7��a��q+Oz�?�^儍�d]� �,��k&:��sh�33�9��.#++�ŉ�j�D^JӈY
���lw�"F�W$���j����3@:���=��p{x;��|>��� ̾�%T�pPh�"�%��Ƃ%�6��z�W5��Ѽ� �Ɵkh���ɥ���}���>���\u��IA���d^fiD���w���]��9^%,_�=���z������E|�e�QK��F����1%E�l�>��^�[�K2��{�1��veq�'A�E�M�F�Y����e���r��D�W`�ѻ�y�z�+I�-�������F���;-��uA����J�r{�D!�t���v�kͦL�Z/_^gu���+�j�}�����[�1��ߕR$�=7�o��'��m��H�y�K���>��>9�&m�
;ԑk:!����2�X��Z�aU����/^\+T%�?���b[1�#�\*�cc�	P䵍��`�PS�j6��(ߣa �p�
pyUͶU˔ˣ%�C��	 y����z2�+Țm���gK��p�p��
�ˀLw۔|��	X�����*���~���pd��uP��V;�q�w�� �!�z�nF�Ʋ욅��(������ �7�t|$Yw�1��i���'�io>%eÕ|8f�O���wK�Ôs�v'��u��a[d@�O/��1�{�8�;u�0F�(6WVl�� �.�����#�)T��nJ�*�L{G�侷��Z����`P�4�Qi*ݗ���l�@n�~�!kx �<J8��7w�bR|�������7���3��V:g�߃5f[�P�z�:VMs�4�RC%͞��{�hg���H��>�����5�Ǐ�0u �tpV��BO2�{n �o���!8E��a��V4�q�J�"H�j�����i�{C�wtQ$�<�<�t��0�O�mG�U��n�z`_&���^&mj*]g�C@�9�[e?t�\{�Ց�a4����)�ѝq�,y���33������l��?_��v�� 4n��_õQ�>!t��� U4���+J����c B$�;>((�}gܭ,���l�k���CӨp..�p�d���]�sQ=l��� ����Cv��|�ٌ���X��
 \8�dK��'� ��b�4����CUW6J��W��=�H�A�� �?��9 �o��K��1�� ��m�!�n�&�����(?�W9-GEE����WI+��[�����%sr|��̙���W�L�r�J�J�R���Ǘ�o����?��U��$n�"})$Fz�(�$�0��Δ��ЎދŏW�D0+|�IQ5��5�&<Yr0��de�䯩u--Zu}��yۤ�_�\�?d#J�_�(p����+ O
e��m�|#��	�I���5[CB@/am���mV��X>��^�p}���[o���S���@?w�Дm힩>/�91�4�NH�� ,b�bA���mfFr;�آ������ uN:��v��a����7-拾�>��A���)�{�Æ��)jW��޿h(o���`�$,����C'�ik�v>l{���@�PXk(���΁(�Y��-�3��>�3_��p�t��]�F�U�C͊��W �.���%J]Os�����^��t�䑅���d���܌�����5ˌ��lZP'G+��Ή@)CFl�T���{G&!�{�ebI���=����9�)��@��9�E�-�/*T��=�1Tp����:�"ע=�C�����,��q��D`Q����V���@kF>`����l�J�]@D�z��	 ��{��bSo��]�����ߤ�9�����!�����+ �g����Z��q��I���ep6p i����@L���#�Rn������tЉ�G`�3�\���ހ6
_���~a&�!M���D����Ơ��8�N��0�����.�����A�X����(E 9;��0*��}�� �RRK���{��v���-d$��[��S$��F���X�3���caa����qL��Q�%W����̉k��ګ(�e֒��Q�Y�|�������亐�� x9j1��y�;��� 
�b���EJ�)
�؞�;I����aT��`-�䐅L�f�#p3� I�؀1�G��'|��U��W�ď��/oT�yKl����c]+ ڀag�5���2�j6�MR��b+ �`�Z��!b�u�}:��Nr0T�����l�U�'�e  ��Ol��(�mA�@W�"\~P��w��4���}�e>�2�V��Z�U4�>c�ľ��{Q��c��J5< b�H;�M�E�OJc�H�ev�ah�����r0�|����`�9(1���5��!bU�s��:W�����+X�H�l�ʊ�����;��;c���?��M�N|消������U8�ۖU���:���wUӲ���L�gaI�W23�eL=k�@���{�l���^�Vq,QZ
0�G�iD1s�h=����0������}���� �3��=&�y�x������vh�m�yQV��d�<�h}�#�\��,/ ���q��S��/K*����)���u��1�	�Q�iC�-[�������I{$T��b���ݢf�u�@�b��/��=`��)�.'�i�z{踎�؎W�)��C5u����˗/B�6�(��j��EǕ T���+$��A� ǼY�����T�p �^0P4fEc)𪂀5
��K D�:�0'Y�[A��+/��Bf�ļ�f��\����S��a,��D�n\���P�����lߓ�j�o���x�Oy�:8�f�;A�2��/�o�5gm^��X��K�z�aΣ-�_(��fz'�ƙ!��yG&P�<���
׹-�Ry�e��mwު��s�x�E��.�M/	���L�6����歱�)�(T���oq ����cQG�vk���y��|�Jɉ�����X!�Vz�XDg�X��k��&�s�Am��icX����pT�-�����w��j�w%B���OK��/44b�<���H6=P�PL��4���x���h�E:�:y�99!)Ǜ)���0'=���	�m,+�/��=�&A)������O�n�+�UTK|���V�3� ��ƞ�#J���f�V�|0k0��gm����O�;�/�IJ��d��^ R#t�
y�r4�A��O���R�����d�_��xZ8�[V�)q(�	dj��$�������0��漓��~z����bQ�/�Isu~w��}�`w!5��Y�����z1���ig&B�hڈ��	�^���\~�H�e��!A�	��⛿݁����N AN�q��qT�^o��
�H�q�1��Q.[�!��O�A��ra��P�eќ��{:�L��f��͕T�Q�;c��=<=���CX�5�g����9#XN����΄���թ^�a�\�P㬺8���۽2L�}��n�Un=ןS�k\)w3;�P�(,��涠���)�9�m�C� ��"~�7��f���\�!@�� Lֲ��X{"�r4��mF����'H쯽�x�;��4m�F�X��2�a��mx	�IGqP���ץX�eL����	�	����#������'�����$[³���=���ni�M�ނ5�.�w0�>9�l�������jⱄ7�YV��&�7�b��L�d�޻}.x�hj�݁,��>�&�������/��U��$Lb/3h���b@zTX_��_լ�$n�eq���u��h��=�Z�zz���f������84�fAY����?2�z� 3�mu��\�G.�\cQ́{����g9`��M���iS?��G��^%��?c��0����\IZZ��������'
��M�t��n�#��
n�Qĸ��H���3�*���?��9G?$� P*���RH��e==��(�T��6 �� x��8a��F&]'��K��G���<O��TK]S�FIb�8*�@�/}��� DYױ��C�(7���w�0I���Clk@`�@��M����?[=��rN�	�1+����l3��[Wq^u����o�����?�P��%y��)�x��b��GL%׊�N�]-O'��(-F/ޣ4��ƍ�^ǙVV�̢�フ��"qo<��z���f��P������&u��N����/�o6J���|���o_��VQ7�}:�����3{!.R>-�>�.�k�x�ȴ+k}�3AEO�1\��=�vV��Ee�'�J��2Ӫ2l
�t��n
��ٮ�Z����2�IK]'��2;&�D�'s['���)���-��_�6�+~'^Q�"qֻw���TZ�xvt��5�Ʒ.��:0D Hr�~';~�H�_ŀ����J�z�Ks���č[\cqn�J!�^�#ft��^�5��͘|,0jy7���`'|�mR|��Ç��g:�s�����1��%��dOKE2��� ���C�XP���q��tG���ܹsqCs�E�����ކ*��-[�$ 3œ��ŵ�~z���)��ǎ��oF���vY�>��Sp|01���j�hȉ�k{�Ӎ;&:����xc��y��/b^Iv��ђ�ʪ,D��t���+8���鳋`�����8t8�s�q nLC ��1�T��J�B0�bj���M��`���o�hġ��jDL{��Z,��F�-��Bv�bj#[,����VJ�$�n�F9�'7&_�t:A�N�%�n�!�94n��
��$��\!�O�q�`��Fg'N��s\��޳G+K�e���QRZ�����q".�b����-�R��V����*%�e�.~��h�	X�`�������l�
m��s�73fecæ���1o���6��fc{̮�T(Qa^�a��닰�6WEycAl���.��tn�k��-���,�ʬ%%es��T����8�g!���hL��e�y#M�{h��m����SA����o�$Q��b��yC%�,,)ގ���G�cP[�J �0¶O"c�H'1Ţ-�	�-/����`9涪�K���\/#f��u۹n+qh��o�p��+4���-"����eP�5��T�7=j��ԭ4�0�[��}�a�	X�DI����A+�2>h��A�d{wu'�����$z麍S��k����1��uv����i3& �2 �������c���;>��!2&f�;47����*[�q``�M�G���̡N��N�#��>�� :��آ��
�ͨ�P��)�h��U��Kȇ��K�V�Q������ o.l�B�ꑼ��q�$Re�À96I~X��2L>��1m�vu~�}ؗ������Ne��s�4��Dugˌ�D��ac@�RaO�$Hm�_�/�z�� '}��"�M���\L�cm��@���_���0��j������}���~�]�m�yɓ�"��pnx�d_�~��2��Û�M	P���)~d�
���ceT��)p!���\�2J�tӮ��sP�__�y�Y11v�[� ��\'����"�Fp��t�-CL�L���{��t�3ɤ��a�X���˒`W�/��U'Y0��g���,�������*c���B�����V���h�p=������K�]"�-��9���=S��\�%5�����{Z��Y���Z���|�m2�H�#)����Ͻf����6k�d�ٙ^BAA+��n_Ox<�g��r�����ZK��j>��n��4�d6��V��KB�H�a�Y@Е����@ܐ�Z�~l+:�2+�7���6t����h����׭r��2�ܛ�t	�0�|���;�S�_;����� ��\���~�7x܍�����D̅�	�����`G|-_�}�<�RF<�yq�u��$ʏ���?���&:ם�0(�y |������ /��V��x͚%�T�h�惭Gv���g-ꃉ�N��e��5�W=��H9�����*>��yX7;�#j<	��/ҁ��f�\L�VG�A��[d�����<�1����l���3gs�Y�GO52심Ȣ�Ä)���n�$�����2yBC�in�mΕ��j�{�b7&v&�tѝ󢼃{)���y�I��Nܾ�dJ�w@D����+ͨ�e�a2q$�����?�3S��O"���R}���$���[5e��vdؤ�����[�d׭,�B.7A)@���$����E�F�V4��F'P4���U�zɮ]��H[��>0+:�����dê0��.���>�e��'��}��v����q�F���tF��h����T�Ql�^)Ly4�J������R�΄�f���^�\:�z��a�~'�T�a�^Z0�F	�Oj\��jY�N}j�r�����)���-&�M�7"9�U��l�t�=A�</�=��Pk=�^����"I�=�L :����+�0B�C�����{�AB/t߉���I~�j����=)���p��N�({�a��ˉ�W������/۴+�@<~շ h��w����.0��"#u�AW0ç
����,k���vni�\�b�W����"(��b>�IqN�	6�S�P�~�8��.d�vf����3��/�1��Ѫj��	��W��ؔX~l�K� �V�y��2!�ȗx�0�Y����@.s�ϑ��\��Zk�?X���<�l�ݢF�oέXŸ�I5�x�ٲ�{�y��r�׊9���;�d$� I�塀��z��q0 6�Fx7r�s���P��H��m-�h���v�1"�\�_��R:ቃ����p|�!�L�O�l��թ�T��(G�q\$��PM�+I�*I�Qr���`�7:y���������֦�%�Y!k�[�.[��z�j��a٦��5ca%��9M2��UB�j(q6;a:@J�"�b"5Ppl��&�F�!�@�л����S�� ���N�g�Ė�݇p�f��9΅jaw���Lre��lNxwg���|�d��g=��Fm����lEGF6��D{V�,[b�E(nx	*�^�@H�8/|�[�s���j�r��r��V�q����{�����R���ħo+�s�m�I�g'�r������Y�\��ӊa�[�K���Ŭlء<�gO�(�鹽D�����er��RM�	q����O��2V�7����TaK�e��ZG@t
��n������v�!�\F�+qC4j����j�a�?��ڀ�RP"�I���V�J��'{=�{�sNg�v�ߧ�ʡ!<O�Jї^�,�+[y��p-���';K<��Ks%��+y��`�"��nYQ��vn	Nz;y�͟[��Jv�<��!�l(��,X��	���W�Ȧ�ʩ����,��7S}k:�!3F�Q6����C��9��B m��e��*��_O;N`C�v��q����щ@���8��N<���i�|�p�$5, ����e���#Ř��hITu��H�X{��E�z�bO�U���'8�3�۰ɾ�ϸF�� �Ŧ͕IIt���>�d	�$yDJ��)2w���g��ˢԩ��2 �ۋ��z�\���E\�`���H+/�~����$ cڞ�p!�-���� xl�`��2�\�����6e��n�3#��tEbd'���ד�^���N�[�~�n}"
�Z�l~�����D�ns@vx+*Nꆏ��@��u��Pj[��u��H@{�2�Ј�؀��4 �6jV@~8:�(x4�C��Y��}w���˦$%�Eǋ�����5"�	��r,=��	�H�����҃��3;`���40���?sJ"B|�yF<q���1�罹������l@$���=�W�Ӈ�-�H���b���J8X�C�Ƨ ʾ[��~?$��L�?���0i�q��;O-�OG�6���]��7��\���'P�@w���-�AT ,:��Y���q��u+�ᠣI��5f� �
u���aqd��dq�(��GQW����L"v�"OZnͷ��[�D��L����/�~}��e�q׸EX��Eey�++�I���v]=m���8�?ߟ���j�J�� Z 7}�]C`�
N�����ϳ�nM&aG�<�B��Lk��TGvNջI��.ѥ9nt	���Rm�&O������|O��U�E?3l�nqh�Ϋ���ɭߟ���|�)��%�����V��P���z�h=���)�� AT�銞'c���WZ�Y̬u@<��
Dc+CiO�� g��/�h��p���p:��m|�4�洐KR�p)l߮@���Gv��_-�ҫ���K� .�ޒ	����c��b#�����aG�����|_�MS�+E7F�
�)~�T�1��gEŮ�N��,a����uyva�����5q�U�}���O��y{�E�ӻ��Eϒ����N`I�Ȭ6GaOz 4ůq�IXk�p	�%bUu�(+_�(��թ6�y�N�����xr��Q����@� �Y���'���Jt��}�Qb�.����<h/�K�`����UK�BK�<h@uc��u���CG�������qqp���I�s�NZ������Xx��(���-����*n��}�,ѸI�����@���՟^�5�ha�~0����l��������+��JmRA� ]Vl���6�R�W�%���ԩ�^��9X�S��5u��ݓ"�z=�@x i���Ufy'���T��dU�<s�px)���U(�|�.�㵽4 �ok��V�v �´���L[���&��s�qQ�w�'z* �1^�~8�
����R`�z�S�O5�C���7�`y��d���/mJG��k�*W��y�#޴'zU�(��Ks� �n�!B���8 ����aG��&8"���ew|ŗ
�ؠَ�Z[ ��K0�Rs>�11����U�j̊E4�a����a����uxq���{s K=@:y��Hl����F�N$�i	�U����=��Y �6U�$�N��)~�oD��\�a�e�;1 89� ����������c��»t$�wWa1�R_o�y�rMj��� r�GJl�c�����r]4_�oix���F�<����g�h)�#�>�̶��98�`\�2+h֝���yR�]Y��ˣ'�u�É���p	��,��0�z����l�5���.**{[�0�����(T��Z^
�88��	���r0K�.oh���ˁ���x��ڶ&@R�<`��NF���[�mC�Ҳ��"��s���'������������w�ѽMWH0��w/�cc�"�n�>^Q<kQb�#Ⱦ��3���<D5p��1����]h�紟b+y<@���!�y6��_��v{��\���{�11G�Eo�nU#C�~r/��|7�+�c�%���\�B����ď6�+�ZT|���<;��U����k*kۆ��:c�6������(M��4�c("]J�'C�D�5H�E"]@z��[ ���k1������~��w������k����:ϫ���x�8�������jwg`ٝ%>�M3��&��UvW {���o�\��U�ܖ~��&qs�t H��9ڂh	�lۄE3r&Z�bۖ�>��,��8C�	�����S��d���6Sh����I��y%��l$�F�[�乎��|F�8��\��V1�8�����K�aĢ]�aN���9ģK"<U4�쨼�!��4�b�i8��<�:���2��X(8A�C�\�����)'�B�<� G�"6���QK�֘F.��������� �X�AA�2w���h�o�~ֶrXq'�-$�_���m���mQ�P��c#cE�1o�t �-,֙��nK1�*f�b�P�2�vO[�=^�6X��I���BV,�y{��""�����g�2����x��];��m��;��zkW?���ëd��ހeKG�=`��z?� ��)Ͱ�EX�'�=�;98+L.Aݚ^_ ��[{%���� N4.�2@^�b�����+��m ��c���n}r	�o%;� &�%y��s��L���1�a���u�?���[k`83@vK�q�$V!���:�I�� ����b֣pY�e$��=�Zh����	�����H;���*_����7���͇���!�2�<4{�Q������k i�X���c.��Ce�
W�+tQoC�iN�����N+]%�r�ŏ����[��*B��F�nȼֲ;��#pWMG
U�/8�)��)u��Ebu&��M�`��pߝ��.n[[�����1��UG�v�������΍��'H�(sDD�A����:��K�.�]�K�.b`j�ur��7�b&⽴h���陙�{�+��f3�t�ī@l8F�"ʀ�������_Ϯ��nº^X/b- k>!|��^�����@�M!o����(:�>1פowFgw1���Qy��ab�눊��Ɛ��ƧZe_h�`�;j1V���9��f�C��s�ḃN��u^�t	"��\u|�i������?��� *X��60Kl2�D�mó\G�a�`98�B!�<�Xa���j�v!���[L�.�>R�����̟�5�ﭱ�Cn+��|XYߔ�����wiN�:θ��-�P~������Uʵ��F)�b��%� ۬�sN�+'��l����`�K�s�������+S
̄���mz��h1{���,}pGAA!��Uf1��I��O|Do�j>�p֘(�XZ�a���V��Y.����Lr6�`��P0��Hq�Q����&0�C���L�/�{���!2d�J���k�͚�{�$��G`����N}��<���N�2�߭�����,�GͰ2��Z�`�D����k�Úù�����$ ?x������֌K'�ka��z'== �0)P��J�������O�.�5`��m�<�'����ŏ9ŅU�Ȫ�ւn}���`��Ir�r'�O���b�T�b�>�k��&e񯴍D�QԖ���_tz��4��0���'�Rb4 '?�"��~H���L�����_��cx��q��ڏ�h�!��ĺ�0I(Q����l�ݵ��-<�V�k�����_k�%�j��Q��jB� <���}XX1�L�,9O��Аd��\I�5:��1�*e�ڱY2���|j��I 2ZD��3p"�ψrB?c��"�,�r(]��@���j$ ���J�=������j��@Xܣ�(YR����ۜ{��%Mp/������I�В��� 3۔CX�	���c�j�%���.���nN�be��eV���c��.�x�"���;W��uY���Z9܇�F���+��݄5!�S^9���(��t�e�^-d�OGh	��T8���Ȥ�:pf���-.��|E��~!2X�Q T�l%�����=~
�����_d�ܼŘG98�P�W��N�r���-J��	H��Z���e�^>��;=��{l���t�y�!8�W  �냵H��3bu�+���|NP������P���z��D �)�:sA��D�W�}��wbZ����?!��rtt���izlt)MN��w��@d��h���󼰲��k��=3��?NAH�c�'t� a���K|O�*�`�C��Ĥ#|̓#h~A�&���4�<�
�������X�SrZ)�2@���F�&/�.��y���~��MJX���M���/js������0P���G�Ze�\f�ye��Л�3�-9u�D�r����!m���u���#���X�9;c`A6�L'�V����MSy�	�t
�FwfRD��ΰ:3����9�>�dg��"�7�"�uj~���%��� �-ƌ�aK#�Cuh����X]+�6��;q��O��@�*1R�>�ѣ�i(����\��"j�Grs��N�^뎹h��J:���E`qݚ���^��߹�9�@�3���1"���g}��8߸&4Lg�:�ڗ��� j1���&�8�����s���O�y�	HJ��2�qQ���ɽ���.#�2��lv��.t���'��P^m�wi~������-`M`�F?0�gq�[���+�Y��$�J톏�Dvb���r՗ޣ�k8�mL��~��cX<T�)�?U�
L�i�/T�����s�ц�F1��b�+Vj���R<�`��rI�P�%FF,���.��J���Jf� 0��\�\�{T��G��{~��[-Z��밈6J����+���8�ypGk��ۓ�PV�ž��O+<��?o3 Dk:�]w2Z_��=wy�!��o�r�q	_E
<q���L��'���laU@A�c��y���W9봈�ǁ`������W�$�㔝|�f���K���z��2�ݤޞ2z��ţB�=�y�\	$d���X��n*(o �*d3$].��ؾ'����8�Qp�`������]�6rՇ@�����1ӏ;��;M���	�J�\��L�h�M`��G�ze�"�v��ڽ�A˶�c.'u� 홌�R�!�~�fj?�,0b���b<�߁�_��!�O�FS� �X�|Y�m-S�F�r����1���&��]c`{��6_���*-k��D[H:o�Ko��^p�p��Y��B�Bd
(F�~��j23�pH��y/�$�d@t]�h駱�T�T�9khh���w�/U-*�H���
	ƌLF_�7�|��Y��틙q�vWav�*Ƀ�2N�GÚ}��E���}憸�p��y����ef���ݯ��e)�8�kk� �;y�C��;�S~�R8��� &��)d"��{�pȭ5>�vD��͆�ortl�k�0����t�7rq��0D��>�9eEJ.�(�N{���,-.<@9���>������羀sr����G� �0l;e>�3�@a��H���H? ɽ��Y�̉P���2�x��3	�
{��Ո�Zȝ=�#i�Of*Z �'	���)�����L�)k����&f�ZJ�{l|u�Y.X"��#x�F�2��[e��.�a�
ۄ/]�lH��>!�e��h��ڮ�gy�?`�m|���E��gp����( >(R�[��'�Al-�pʹ�Z<�~��6R��q�}��s���Rw>�V�ژ��P�����U�	��"pC�&�Hlh����n��}�@��,�]��3�t�q���N�yZ@0vr�yJ��&��h�ס�?x?K��6y��<�-��� *=Ȣ,��L��J�U�za#�U�nʓCؒȨkH��8��W&���?V}jcX[���0M�ټ�1�ƚ�`c$�̼̦��|�=L4�
�%H�� US��k�\J��_1��1�r�<`�"���9����]V����x�-���`��#~�v���_���	�\p�����aU0����2�#°:�%�`�p�E(����,����9i�ΦB�^���u%+U�(bXb�Q�U\~:����a6��s�c`�(�����04d�v���A�p*-�Ob
 �o������b��k�U����C`;���<x��'���.�&V��toᘏ������;��Ҕ�I�M����;��)&�����b��$NvMז�r�:48�X$�)�	�Ɔ�?w��?��7'ϙ�����3�������a���(�u��Q7l�:R����V���ZX�b\�A��+���ɭNy-�>,H�SC�L �� k�$`
�����-�Bl7�� ��Ú��rw���O�π��U5�b�,_M``�)Vf��S�]�+�p$���l�k){�pfp�"GO#�sC��"6�n�!ۿG; �t�/�+@j���3��G���B�m_�;�2��/A�&��Mp"62������|������]7Nf�Q��+����`��'eQX�� X,	ڙ�C�.G4�
yĩSǕ�Ѵj�����<C�U'~�1��'۷?=���(j�B��Sl��z�)c�6|�9W*�1H�OXI]+���M� ,'��7��e�1���@��X��;=}�CC�d�@�?�=c �[�o���*E���������V�Y�gR[��H[X'tf�"�݅�ܰCg����u��(�*)���N�ߏݧ|d�
8���\W�A�sF�yx~��������#Hh8���m�����l������:o70X/��$]Qh�j�%��1��q4zm�!·��SO������z��[�84�܂��|�F���X���q@֩�����g�[#nia�|O�E��a�7�γ��6��n�
s�ziH%��D ���*��0X��#��a��R��p��o���9zs
��9ߍa �Nf���t��o�3k"�`�z�<�=�_m��X�X��;���\��aE�i���R4���
88��Jۘ��x&��:M��lZ�gM���9E���Â>��(�Z�Rɸ�%+A��������̀y��_]��enQG �c��!�1��yuA�pSN���\��`�	������P�5����hy�Y��#�z�T�e<�,�2�Sÿ\jE�[;*�;���������M�?���~�;���}4(���� $���;�����.;��tM�E��x�n"��e�f 5��S�|+���Ӏ^��~s�_��+`h��$a=����*!W�LH��c�d�_��@��6���b̔�� �6R����2���y�m3���՗�FЅ����������ћ*��͞0**/��,��!���e�O�_a2��v��7U�]���-����@��yL��GҠ=� �p-y-���Zf�w�\NX� � ��w��4�&p2�FpI�-�m��n�+�+\��D�$Xeܺ p����7&�`r��i��O���,��
ݴ/�x'��M.�{� ЛF𸑋�볝X��$ؼ_#�F@k��轵V�3#�M�� � Х��%�5�eK@Aϩ K�V`�8p���Ɋ�ڑ)�+�YE��m���K��Kk�Z�w���t�r�/��E�U �]����/ ������l
�WД�9QģM휭".a;U��7f˟��=���_���ؕB�j���T�y"b�?3��ʌ`�K,ߓ�
��0�J��s���� �	��0�0�B���b{��Q���_f���)�Y	`"��x-�<p��K`� ٌ0mxӭ-�~1���:pnL����~<+t��c�Z�����0�9IG�D�������F.�fM�=��>m�Ɠ��cN�K��V��|��Z�.q��Z��+���S�H|kT�������7SA�W�x�W����!�ϛG�����������'7~}q
����O��"��������;�2���{�}�ؿ��;����:7��Z��{f�� ��� ��� ��A�+Z��{��z����Ѣ�h�\NoՉ��|������;���fp�����w����Pq5���*��)J��M��x�hw��$�0�al�.ŵ$u��4�?��z[O]F�pB]Z]��y9�?�v?�h'Y��V����T'��Gg��?&�,k��9c�Q�딿�v�?�F���T�M�g�������K�������_�K<�pn��;m��1.�	cC�����ɣo�pX �ރ������ٷ��l�?����)�&�ʭ��u.�"+��47����QL�:��K��Kl���v���p\��0�xi�����J���>��_ߝefb�P��I1��	�	D<��VƂ8�DI���gɭ�j}�z���� �'�kg7�/[.]���w�:p����QT�<c�i��gR���C���Ks+����%���UJ��B��ϑ�ck7����T�-��U��0�9��(?~���X��14�X����#�s�}�	���5+|��m�t��Je��޷�0����Eϲ۝�r�}���e|��o���VT�E��F��b!��4����`%N!+%M�����@��1�t���a��n{5y�+��1�Gl8y���븡��������\?XϐMe����������K��$���/N�71 wK�*�G��oq�>,|�
Y�#0�`�|P��S���JE��?]�J��h��y�������(Lɶ@��Y�zH���˃Aa��^]�'���*5C �%yMa2�Ky��b�������(��G?����ݙ$��`Gl/�m.u��N�F{�%�Ā�x��oC��p���W��1�AX)yx�������f,���Uʁ������c�@�nY|�N������Vן�==��ү��p�Ji���XOW��(���ᢥh�_98��(�$����]����������H���<	���6�S��w�K+�0���.��x�,D��w�����$�J#�{��"���/�����%{Xm��_�5k��G����5�BV���[���/�o�к����*B�܌m\�g8����̮!ti@���nR���|��\�Ա �%B�E&���o��e�}N�Bl�7��p�熰>'7Sv����iJHhH<x�~m���A�Z9G ��G��[a�#|��pST�e.���^��o��� �A���)����M9 .���j՝�"|�C1����o���BŻo�������Y%�޹#�|��͓��	5ю[�F�0�Ho !�nBм�N�A��1i�x�����`��E�j���!&���ウ�����~#�g�#� 6����B��^X��&�0?%�kss+������Ռ|_\�k�r2�$QA�<�x��*�h���HHN-�� .��&��y���>���^��z��t)>��#~\�b�~�����d.u!m>A\����n*��n�<�sՈ�R�{t<�9	Ac�����@\����S�C@SΘ�*�ط0bf�p���(����H�^��}��ʅp}=w���W�е8W��t#uE�$������}�r�M�`S_jc���[��A\ȀC�x<��H/���c�����@��\I��/�!L�:���1H�I%��ʛ)[}�B�N
ڻ?P����Y��<���2lbF^_��8���͟���w����ó�'n
:o_�|��4�%z!�og�̊��zUO�^���~��Vwd} ?PV�Qየ��~�/�)]��Z��٧�	Ǉ�����8��%wg��⅐V���_C���&[L�ݗ����$Z�Dy]	���m�e�LV�;�(Ɔ��+��,l�Vڄ���p36�&V�B"+F&K�R=;������ަ���f�[3�J�}}�w͈�r,�\<��� �a��D}�D�-�~�1�n�ӗ��{u���ܵ���Mbc�������/9>��"�����"rAp՞gi7�pR�H��N��V�Wďg�f�+D�h\���AkE̼V0���d�Ob�TE�@ЊϠy3o�c�2?{�����A�i�Up]'-��D35����6�Q�=v����c�ͤ�3���1Wũ��嫥a3gR�'6dk�/�ٴ��H�|�I/��R~h��r!�8�7Z���/��)�+|�p���h|��&,�̆� =�Ւ��\7΄p����M������w��{`0;O��w��㔜|�U��(�yɥu�a9z-�y1g��r�����̲��]��HYv8���S�:ب���^�Qj1tk]�[zH00���R���uw���!�Bˏ�����J�cNh�U���Y)��;�AlH`��2*����=E��ʹ�ͺώ��?G��E)��y�u�K��OϤ#�S����>3�/���M���0�k��(?,�a-5`f��ER���Lw(�`���,b�	��Z�L����l�>̪OK��d��x�b�����c �N�J��W$yO��а�vp��%�����? ���k5E5z�Ȋ��{���I��n5܏��#X�N�Yv���ݘ�!w��b�c�l���K���OT��x�����3�MS]��i�&���q����R-�x�9����ӢA`"��	siCr��}ˬ��]�t+��G_e�m���,����$�q_;�W�\��W��}<r}�*WxsjU!�tq!p��/&��J�;��������CU1'2�����g]��_�6B\^/0���['�*}��~�+��������)��`/,�`2{��_��w-�N!��	e��_L �=���D�a�ѰeĽ��i����ex�2EQ��
�NL3�()�j����S� ;Fe���PjkE�x5�L�.��#�f_�^���<eĿ�u�,T +}lt����[3��$[?��!p�Yg������i����;�K�!��WI%���"�6>��D-�Aԓ��B ~4�=G��;����<�4f
�0�W�p�Kmq�^}:)�h"�|Qek=���d#z��6����a7�j��FL��RL��h�!���q�����9<��Rjb��c�^!z}�ab�!���'�ᬏ�F�O��_���˾�&[9Q�;�QT5s����,� �͵x�5]�_�ƝFx[6��PNd�߶�:�8OO�_��- �k}}*X2��V�a���h������Μ��W��-�~F|�'�����K�|�o�[��ڔ!�F>h1�DY�����������t��5��X�w�R�HB5qY�{7��O�_q��M�Ե �|V((^yx<l�<��ʑ_^c,e�G���".�p��J�G.����t=�x�}4�O'/�\ꄨ��Ұ�X�$:9�x��#8�]��e��㿿on?�/�U	��m���慉�'�m�)�;+:�j`��G����e�!�y45�X�7h*s�R/�i�ǡ��N9����⃿2���밵B���h�t۰9,��F�{�ֹ�><\`����&GsQ�s���?N���B�J��%��9�i����}���\�!����,J�$��1x뗱�<�z����r���".��k}��>?��v��Y��$�vᬊ��;�*����f�#o�65���o�B�A��v�妰����}��CL���x�q��'��|ƥ��54.3<h�ٟxY-���B�A&?����k��D�k'Nu�X�;K2$����{���L�l�F�2�7�c�����RJ����4���9�@��?��h:ǋ��<�a�����)Jٯ�Y���Hw�C
���zQ����wEjq��l�W�8�G����g)%�K�"�P��X-A����Z�� C��֟k1"�[=W�KJR���*��6M23O�n�+0o���Y!�x��q��R����c���q��6����_���*J"�΍��W����J'���:�9����HJ8n��35i��������td��~���ʉ��;H[%>�X���;K�]�bF{٪��Α��z3��G�?���j	
�=4�v��zƹaN]y�q���A����=9���C]��IL�y#�n|ìn�ˉ�w(�#+7�N��Р��ب��|E@<��?N��à�ҧHzV��r�ݱ��nV�a\)���3��B��7��lU���5��N�J�B�M��U��H~�"�Km���e����&
F	oNU�V� R�@�=������3�����N�\�lqM���$�o�U3L�ڶ�r+���E+E}�(�E�]�`9#�_�bC+]tCi^���_+vi�H��h��0��>a_��_���	d�qh�4�T�����Qr��}�Ɂ��s����Q���oI\!#	چw���o�+)ثQ����W9x6�~�*h1Y*oF�J�D�c�.yf6[f$)�,^�~Q�a,30��Tlj��U���0� oGP���E��MW=<�����cg��t������56~e�"�q��@A�}�]i'��o�U����%o)s5�v"o*j_�j��UY�Y
�Qe-���x2\�dCS����Ǵ�Xm��K�
.�>gy��_�;MͰ,��l��j��S��3�ޯ�O$ݜ|�H�2�E��Ȑ�h��p����HD���D����%Y�y��1�yL�K�y�u�A1��!.L��7���Gl!l<*:��VTt���/�+�J,�µl��#��ݟ��/�m�_��Nta
	�|`%+��#ŀ*]�DE���}���������4����zh۴��\r�"����6T�7E�wf�����K�C�I޶�:�E����73�ST�\��2#g������*]M�l�f�*��t�TH@����h�2��N0rQnI�P�E�U.���ή��|�����#r��]Е�l�����̥�\��㥀F��/���y)+M�老B|8c��x0��H)�����܏�#���%[b��x?�sV;����z�g�On��2P��Iz�����R��K���Z&u�ee������������6yV9�zG��N���45��q�����9`Y�;_fv�y[��5�9�ޖK�夒bI��ߴ.W�Ė�u�\�;vڻYɫ{�������Ո�����
HvWt9320��Q�	T�L/ ��o��v<����vo1��K����xpt�6���>�xl;9ɐ���o���}�¶}�h�t�c�hF熁�C�lg�6c���J��LQ��������#�c g�����V��l��e�2Jn�G4��_+(���쇎�)шA�P\2	��?�3��Y����\���2E�Wh�<�E�+��G�����J�d���!6jV�K�7��W+�fOv�t.��l)�>Pӑwq�*!����r�8����ɉ�؎�C�ݮ��Áfn(�%;��ʙki6��ua�f�������pN@�-�:���/��Rɋ縊���2^�(t��H֮u���NJ:�k)���#��b��%��S&�!֔%�ݘ�-X�{��'�xwTǁ{a�����s�>&�Λ'�|���=&'U;Y�����k�Fz���L:�t���/��,X�bjw7.�%v��ؑ���W(���ـ�7=����u�V^k�Qx೒�a�۟����[�"7/?8$d���O�pSd�Nt0��D�?����C���6�ǫS8D���=����ﮐg��$���l���M�v+���K٬�Cn�g�`b{��־y�F�PL$�UC��;�g^�.����_�Z�4���خ6�4��9�8:	Й�8��֖e��[�l��N.��+"��`��؆YM(�{��͘95dM�C��?����p���J��rN�ZlI55�=.|��)='���vW±�Dʤw��,>T8V���n�2��X����%����?�^��z�:�:�v��Q��N���H���3��۶A�(צ��aSC�N�1�K�CA��_&k��L�{&t�q�-Z���&^w�?4��t�D;�aW(���X7�2���I<�)'�����{w��m�:�K���nf�Q��)�j�a3wG�0G�ƭ�n��NJ�����%Ȋ.h�n�;%��[i�]�h@����c}�p�")��� ��;c�fƽ>�-5䉕�`$�/ˮ�|���n�X%�Z����W����8�Iu�bm����^y��^� ]�g��C�^Q�9*_��g�dF��(����@S��v�����g/N��)�%��Bl��v����*���Ó#.���4?�Z�*�#��F3w�F3���b��iCP&7�e�fb��� mʼ7����ư,��eh��t��ͶѭU��O�~R�6�s�Y�ֳ�<��?�9�2�5��2'l1�jKW�p��\+]B�eoK0��Od�ޙPl��O�,G�c�e�/��Ǧv� �@��5	���S���X�c�P G�ek��c�j��I-v�m:��1Y����ڻ�dy.��HD�#��6��1�I]������5���l͌��$�J�ͷ�ά�V1KÑ�k_��h�j�}�S���P�Ug�����h����>�;p���
�x�Raw���xO�Rop)�Ŵ�SB7y�R�7�'(����+���^[���s����D~�uB�F��m�CP���#筂t��sT䥋S8}J�_~���.��9r���(��I/�Iv�����;v�h���T'��O�F�I/ ;#\�?���.���N�(Ƙ�{i���-���1�m�}P�������ߔuo�
�E;}_��)��h���>�X�����'�Ǐ��=:��ww��/���Q�U��D��b}ZPZ~}�3�x�|��'�[�t+�㹸��Ѥ@��'��	��*��b��媩R�)E��o<����F��[K��[]\�X%_;�����}�����K�?~�UjV��Ag���[j����*76~\��#Q��O�N��@��p�x��ʡ���?ֽ���\q{�@� �]��S���t%"YUU������P��E%���ϳ�n�?h�N)�޴)�?��� �?.������[��^����]اؓ�(e�@��e���LN�l��~�`��Jr�*o'���;���2�X������K��	9{5�1ja��(*�ե�st�ԝ�E���Βt� /$�@�qF�٥Ě�y���&@@��3�I*\�Dr�F�����(��2�+%g�4�3�����ȥ�;�p+�uB9��011ZMr��6p��S��Q�jR�G�_F0��%��.3]��ͧz� h%!Ӫ���,4��������K���=��:�%���
X5Li��$x��B�:~	��z%<�������Ϝ��=]���":��&]phn6=#jĬ�8k~\�Pv��+a˺Қ���|���|Z֣���_m�\�p�Jr�������N���n,X�=�K?�q�^J ��4�}�j����:I��P*w>�%5#�Yl6�Ƥ��p�ˤ����������׶�:�B)v��+��v�9�u4r ����y��X�+�|c���)���H��R5e�NƢ���3�jצ���׭f�ͩ�����.�߭%7&��{�snD�$VP�`e$��mc��".s�{/���h^���e�q����?aԋ���B�4v�7� ��ѳ�w��L��/���Sov0�0��5�����
T:�8����߀Ȫ>x�E����;�q``1ZHw'^Z�O�����M�g�dK�y�)f�|�#��AR�
'Q�Z#
-�zY�.�㹎w�~p��C-��v��?0k	�R��r��I�yF�C)1������)ل���/'#�45��y�:i�Q���)Y#�N^7�ݱ��n~��A�����b��A�����x�84��u1i�J�<B���p����l���Vg�b�|u�q����.:QX���3�y�@�o`�m�G;����E��@�laME��%��O;�b&�	ڜ�w=��b[S��N��|�w���Z7��S��O��C;�B�8��H&���� ��Q$x�n5�'��ɼ;!��)�lȸقyT��x�HFj��Uo%W���-�1l��Q*��yF���n<�* Փ�"�v_������Z�񭙀��e�ec햜Sڌ�m�0��88��\Mr�4>L+���/2:�]0Mm���	-�{c�Y�+D�o[e2پ']�:�i����d�>�1�æLR4߼
ϓʵnV�����U/���Hs)G�2�s���^uζ3����.q�W���_�0y-Q��ޖ�� 6���a�|��������R��m��"���;�΀S�8�ox�6�Ӝ�����K����� 8YTH���/���fU���ĉ��e��cل-�\��1KB��TY�����1É%b����K�ɔo�Y"7�u�tC���T����1�9����HZݙV�!^�-qi'WӍ�3��]5���6��ԏ�p|-��+7��w�\�e��K��S,v�2�C�;�c[%>���>W���q.N�hmnn��;�X@�^�Q��XM%��Vr����<���Ej��cG
��ܮ�N��c�w�lS4:�R^ ��t��L��e؊jje�w���Mq���p��"f�6��H�H���l˷�d`u��\��WRRPw���of�8�l���m]����/������콬v���0��p��w|<GbD>T��T٫;1-~�A`���b���e�4[�����S8�K�j���P�p����������e;�j.�,vij��m�B��N��m=Y�z�1?�������=_d��K�s�mA%�<t�bvK�nβ;f7���	RMH�U!ѻ���봌Ø��{�c��\�j6�#���a����ŋx�ʠ�/nt1�ӕ�**(8x��9_��t{f�f%țRUUZ*��i5)�&5&��u�7�\gݧ����ց7��x��}L}�x��0p-k:�_�����\~�����em���uXI�nӺl�����^n���&'9_���u:g���V�D+2�����x�s$o1�F���=�y��hL<-�q���l�{<k��9�����~{F�����a�TW��%[�؅��T�
���C�٦�V�s��;r�$2L�<��ߩ�V!QCM�4��)��H{��^1!'�pW��B���l�;?&G�pE��,�Y�9��P�2;�z�G\&O��cg�+?^��160>�#��~M�8=e����� E�|8H9`&���+dG�n9s2�)�-��Q:-�q{e�}���U���8T�T����OLd�T�����r�Ř7����w)�`�ٳt�0��_E�cN-'��p�"f��%x��U}��9���%�ݸ�Ew8�9v�y�"#o�W̗���'r֨"�fW������~F��j�t�yt��䙛V'R�=��aC$�cS�wA�Wҳ����@u����]�����ô���������U��I���M�ǎ���IO{OLv��1�篲v᏾�d��L��Z�!ʷ����A��|�\��� C�X��ѩr�/o:UY�o�*ɯ3�n/��թ�v��8�W|��Ԡh�����`��6{�L�B *W�XnMaR�����P����zcݡ���
�>Wi�޳[�+%��q�ޭ�(^���>Rc�r��r��zF�����@oyxM�R(A�!L/�N�;Y�78�(�UB�]��]/����.M�)c��o�\}�\��.��T5%��d�sY�f���HL��w3D+g+�P���6ؐ��9Y��:">8Ξ�Uz����i~��q2lg�X9�=�{d��KM!%犯|���-'��I^G�!wF*RJ	�V�c���`�r�����Z<wuQ�~N�7�[��!z��6>-�m�����`u�S�`�[�߀o��qw9�I2n��q��K��ݷ�{�U����/n���G�%A����ٽH
�A\�j����kz�҃�M\zJpC��b�r�3�n1��R˱�5�ڎ��G���~��{d�����g%/�MX�2��;��w8�=a�W4C��׎��u�����Ir�	��7ԫ�1wB���|&��[6c��>����>��Uq���u�*���{2��)��C�p,�U���Rc2�c��t����Q�샶rh����;�Ǝ�H�,��o�.�ޘ�<LB_��7+k@��/EJĵl�ꮵ�x�8���b_�ż索q�ݫ5r[��7�?�dh�K�f�̪��R���Uz�e����k����`��ݎ{���������Fz���t��Z7�]�M��~ɿr����'��yˡE3�~$�d�]~5;��ԏ�$��Ão���[՜��ڞy&�+n/�)s\7�:}�F�(zǺ�v ���J����xb�����	�
�Z�2w#[����V���T�ț��5y�I1f:�$a/�j�ƴ�CVc_j�Jw��VEg��C�f���ޫ��}'i<?��¢lCN�������[3��gz���rL��PբW�6��x��6d3ҹ�ᑵs�R�%pn����>�/�2x_k#��;�5]C]�����ǭ��u��E�l��>Ta�֬����?<�pj��*CX�=t��>���S��� l��dU:�il��or�m�d��%������v��*3u�V�����M)bn�)U���מw}��Y�݊р���Z%�������N�%8i�������D���&��6C��J`�֗��*F:\z+��=��aN�`�D�^ٮF�$���l_���&:y��qkb�-�W�4�J0���s�M�]�[T�^V��o`B�N�����6��n2���n��!��6`��z��~oʇ�z�v�0��L�(=�ҿl���9�(�dЏ�|xc��q_�ڣ�P��7�n=�V��zz�g��}��L���� ~��*�`�-m7�\*���2�I|"U99�3��G7:���.5+��ib[����릏h?R�"�&���dj)[��A!Rt�źj�)��ЀG�M$rȮ-vz���<W_�|�;cl>z�#���R���dL*���7z��W�_R���&NVP0*����t"��]�TF`�Zbu,N�y�%67��n�~
e�w�<,��Vɥl¼�H���Rf��LJ���N��&ߐZ`E���2�\���{Diʒ�jE�����wO�z!�{�k�VX�7:�#���j�a�S���P��Џ^��sl5 ��|e�ƞ8�����l�Z���?��^i�xңq�n��ݔ����Zr��;~�1)D}lOK�R�|)!��(L���]����cj8�]����n^4}��r��n���[�0�S@}��|8P�\��.S�4��Sy��K�������%�Η(6,�:��4���q�Ų}�}��Mz*�O?4�s'�1�i�����uz�t���5������l��&(��u��;�� *��z8g������b���E�t��	��&�g(i�O�/�i��
'$�X>B0��.�Wc}�.�P~�`���g�$�v�x�{����n��O��9��ַFq�EL6���nZx�->ö��6��Y<&�Ol�����R�>y)�ψ��)�NoQk�ƆJ�@���tA7���E�_��k�	��r�$���(\ǽH�NT-bC�w��H1P7V��V�u�6���oʠ�ab�7�ո2�!.�Kmp�e^�]s�w���[i14>�w�s;Yk�>��n�K1T�@��pz=z�ϴ�v17�1ì����N��2TqT3},�D<�Ǹ�ʅ2�����Bo,�_�o?�J����î�]�s���  �b̇z85���Z&�����CVo�)��T�-+���l�5�k�l9-Il���۷`f�<�\�=މ��t)%'0�\<M�/�v�]`�����>���+��õٵ��)6%�p�q��υ��j���B璀��|���:���q�FK��1[��t��Wb�($��nq��?1S֭^1��{I[~��[/�ȓ�+�=ѻm����a�..���<U4i'����𔴚(����긨�������Q�K����[��e�nA�C��S���%���w�=7���������u͜9����f������0�M2�"�7�I��g�Ϣ[����-�Ԥ�I��1�������`�h�_~Z"��y�ֹ�J�>ְ(J\�>��4���p�0��lK�J<.���F����/<�q��;���&�K϶|5�����wz]7Cq���1�\��3�|�}��������X'���$��o��|�/�-����>�� 3�ǭ�2��ӯV��,����1̒���i�r�3x���!��w��+�I��ŗ�z�)T��d��f�������*]]s��\D��p���oL! �Ӱzf���#��C�yC���M�S��zN�ٺ�7�(��Si��i��2bB=(G�r�*޷�_Z�
T�������[��������x�D�"tŢ��*�� PX��-c���@@ڧI�&���x���[���\P{�grH�Lzt��[�L�y 3VwɄ�m��[c���zWx_�2���ƳO�;HAee�&�c��+��6ê�����5i���UF׷�\ܾm(�Ҫ���K�אy����Xo��|�>Xx�0����L��z��AZ(Of�Sy}q�Mوi��h$�x�}��hqc�j�(Қ�����3�����=n�~�H�۷q�QΜU���k?����+�ܯ��O�bf�~��v��-_6��a�C�%�{3Dp+�v���A�����-���=���\��{&����1f��l�(�:u�0k���[��E7�)���q� �P��9dQ'N��j���~���WR2�`�Q���T�Ċ��/���G�!�i
N��L� rSk!ܓn	W�u"��vE�'t&�p��7_6};;W���h���~��� �1�~�m�pK�-X�R�.��t���h�]��Q��r��Y��Зr
+����fU�x���$@��������2�s6�;9vO�����O�����1 �E�6��t��W���G��l1�=]�aѧZᨶ��x+{����l�@������f'WIq6QN�a	98�p��F�Ddq�����CE.$�8%�/���\>ކ��&U�W�_*M�sЕ'ۧ]Nîv}����ݾ<
7՜����g8ru� ɢO]�` tE$�݊(;�}T���ӢEzZ��}H?EqF�h�~'��grvC��ڙ�����{y�򴷌釕��1�2�'�-��S��_b�g-��l٘�F�T�.�8�����kW��6�g��,�s�v��|z��7���#���u_*�?��yJJ q�ÎPt�;�,�X�,���VYo�9�ṫ7�7��������
��?eb+'��)�x�|�/�����m}y�z �cX�ī�R���s�	$����U�~�m�:{{���<��ݽǅ��2]�
�}#5F@�s\&��������b��<B�d����x�}_�L9PH��r1����n;
�פ�X_���ד���?��z��YE��Wy	�xk���Z�A��A_���ؗl��\U����g�O�O�v��V4��W���,ζ��PM��o�5���M90I��y{�(co��e��&+ܞ��U�>O�t�+0��ӊ�pwo#�n#Ӣ^��e=~��9�
iu�=/���r_� ce'��[!�H󃬉�����Ʈ�-z�ϙ7Tж�@�� M�-�����̲����)҉k��NT���F�?��6߻Vi�r���A�.����1��뻗P֙�Rd�t�]I��w�ϯNK��C�[|P+�^��A~h��_h�i�wD�ߤ▛yA}�g�B�������Lw��o�F�7۝��#�>f�9���/Rc��������[q密r*SQ��~m#E���O�wф�{ݟQ>}��,�B�"���_8�䶤7��1�DWȔ�e������@*�d̼���R�WDR��#[�v[d��ߓ��oT��k�<�����k�]�D \߿2|пa@��ز�:� {�8���`�c�f��yEð!F-��Vpn�7�����7�ͭ���-1��W�W��_�! {\Z}+����,��Y��V��ߪ��e���Sz[�������~��$���ޕ\�_�fo��J 6��+�ns����YE�����j�-U��� �a�؊Z٘b
vк��Ɣ�^��N��emo"��%�'A�AS�u�_���sH��W�̯�<]�Zg�m~F�}��{r�-��xR�^6�4 :���8���Xr���C*O�������Ү���G�6���v�/�����C�Q��l����Y�}���?%�3ڞ�j3mgv�?˕dc\�����Ryܾ����]�����~ݝk��t�\�E��f�g��
sA!��+˝�A��\��v�<NT2L���:>�"[�hҧ�S6A *��ۺ���+`��h���)�0�o$|N��d��L}�mQ�{8��g�*�R��|7!��e_e�$!#(�]"�Vk�"Fu����CU�k�*ky4�E�{�$w$n&����삆O�����%��M�)_�S��+3{>���vkj}�����L�b���a>��j�j�����<�T�qh޴�lU��ԩ��n�#O+��4;;�oj9�M��䥶d��xagenv��F��M�P;`���.�ű�a�~1�;����/cM�A|�5c�N��$zHkw$l2%���5�'
��G���͞++�fuP0U��[[�����A8J����hĩ���E8)�E�m~ޚ�rb�
�eQ�L���T�_��R��Q�I�'�G�t����Wƥ0��n��_�솱��R�^OÇ�EB�[pη7\AB�|�����s$�˹^T�˟;��'j0%�����T.f����t���w%�Ǘ|���9W^�!�3�i�^q���>�0�iE���83�5G�owf�ٵ���"r	h�^2����H�<޸��v��떕�mڌ��\}|�;�<=�#��j)���u<Hf�\��k�7s ������䵐�Te�_�O�k♢�a`1i��w(K_d�*~1�Z&m�#W���fP�v��do���]����:�HTC=ء��sT�ɶ~�lӛ}�X��Dz�i���/p�s��;N�l��-�u߶f��twp��N�F�j�
¼Р�pd(�R���f��a-P�d��#� ����|�(%6�]�=j�M�)O��C���v�e�CU��d9��=|��
.��|ʎ�����*�Ȧ^�2�����y�"�Q�E�4�̀|��zK��L x����Ff��,-6O�����m�s?���������ec�����E�������ҿ�o$�KG=T�<�.��3s��~�;2R9���l�R�|D,ad����X=89��O��S���$��/���پ]g�.��)�|E�鏡���`(�Dm*V����N��#�`��[���$Q&��R앛�"M����!���p>�P�0*|�E�P.��V
��M-Ǥg$6]��ȼY�s���<� �㕆�����1�.B&L��%\lխ*KCI�q���G�;��,tPG��=!e���苈:��܎����`�T�;	���Z_T�ws-O7�V�~��s9W||������T���Y��pQu)�	�}�"SP����A��}z:ǩ�n�96�/w
����g|E����5��>���߅��hb�zXH�є�w��7��g���
]�F2/�� �����U�e�u�Y�����A��s���s|�MqF������i�%M��;�+��A�d��X���nӬw)�a{�[�n�B����FY�ԑ� :$���My������6�;��ۣ��
�bz����ɲ�U�f�x�Y��8��Q�%�lJTI�+N����/tt���rG�Dy�aԵl2��);M0<-��L�5L���:�iC���rm�����2�����*]�EofK���EU��+�J��";՜��ҳ���uIQɟ4�ғ6�
��b${hxX�a�2m��+y�7�+�c��W�POr�]ì�O����?��IKk��U�5m�l������1��A���9��+^�#4����B�2Zq��s�I�]��/��<J&��g�娰e��q3�.��y����������ը�+��V�Q���e��I��kގ�E��h�	��uZ�Uw$J�"hh���.w��_X�n�.��Г�x���8]gi�ܲ�~+�����Y�0���U��jl�Xx�s$�h�Ե�rT��zv�e¾���}	��w���U�����m��t�~�I�M�&��j�ꄌa8)^��{q�ϴx�������z�Uս#S�s��9p����o�G�	��~o��i��IVJS|�G�8���'-��l���F!�����
D�UW#��	�Ȗ��	��D���x��H���³����0�����Ia����㴳�]��ԋW�d���:A�K�*ީ�Ck���W�8G[�y˱����,���h��V:)�d~C$(m�c)���d8� \x�F�P��1v �����׽򅨁�6��������*��	R���u���v$!��m*����&���wq����T�D��q��y��:z˖�����\$����� ���G.ݼ
�J�p�w��̦\�@_�:)P��xr�B�.��i�a�>ODVe��_����Y�.<\���{�8�&Zf&D"M�ӖK��^
�b��bL�~q-�NN�U�?EQ�q�s%Z��D��{P�0mW�6�#�Ϧ卌��)��W,��7V�������ģ�q$fd��>�1�n�����M)�tR��(�+�mB�>u�i�&�[r�O�O��C�W�t�b$�dBg|�6xK2��ߚ�%���պ��j������9�ӻ����?aK̄��1�ww��#у\����<�(�yM�*m�u�Y8y-	�����4����Ae���~����B$����ײ�AP)�U=1�Ʊ�a���~�}���?�d|`�4�ۭ����ő{c.Us֨�F�$iC��Z~�h�dn�wE�^�����y0s�x����ѯP�+���2��r��R�u-�hKyP=Cj����A����'TN���t�����ހK�z��^��@��`��[�x�����o��Đ�e��[��`XM.�D��ƚg��.�_;?_y�,�q>�V�XB��)S��e�<X�3�[3n������c�1�*�h;�}�!�cJ�yW1���Be���I�=���ؽ����J�DV,�Ş+����|Wl'��7����Z!�SG��y��+�<'�^}�I��%�y(j%O��/�2`��*ݾ*0��F+!v�P'�\����S���~C��dL@�����2�,"�P�)��� ����W8If��TUf��fc렫��=���\�6G�±�_�w��f�'�wl`p�A׏m����Yfr��Dc0ݧ?��}�(�<@��Ejy��@��&o�[Yr�{�������u��x�B��Wd�LZ{$˨z�D�.���xJ1�ZK2�ڌ�^Q��`���b����w��A=]mͷ�_�dz��-��܇�����uJ��߾Q�O)sq�.��,&(/ �ڽ����.�D�b��p�'��B�r�V�"����}���[��U���O[����g���u����#.k�p&(�`W.��� ��s6�?C+/��d��b��r�8�3ײ��a�'���k�	����:Ѕ��hƵ�dCr��Ϳ��a����WJ�J����y�\c݅l>J�*���i�r(U�V��V�����U���Pr�I+׺��VsYr�/⇛�����D<^�	��q�`�{���b+��<����yL�6F�6z��r˸Qf-��)��r HK���r��w��v䅵�/|&O4nH�����J��?�:�4Q��-��m��^E-Hc:�+� �YX%���~�Ƥ��m����E=\�ߝ5cm,_3\-=�s��'�����G-C>�7�@�z+�Gϯ?�BGS$���Xse�k=e����j�9N@�\�x�|�t������ݭ;$�[������_�%�EC'�g�F�bh+�m�G��S@�uR 7�^�K��0� j��͇�3$���B��C���5��ݟ���}۶1��Y��+���5���O�b=.�0-�G�zQ[C����dLm^oc��㱭e�`f�C_�һz6�g���:zf��J��1�A�#dyfp�=߲�>%��>�D�� 3�"J>��Vl+�K�^?𾖌�Ř���@,�$�͈wm�j�< �V �w������\"IN.�l>�����:�oY%�3|����:��_V:_?n)�"����[5@��$����ˑ�c��=����6��0v�:��#M�m����]\����6L���9?l���y�?֚ͅ�M���㉅r�_1푙�!m�6s`6��!?,��������=�k6�&�*����[;���!��g/?�h�z�uH�^z3Pd�
:(n�I#p�ʄ�`��)xe�H��3R�Kg`P����M��m�*�{�a�.����*�biOb~g�5����@������S���b�y�rq�/f�Ǳo@W	%��W�7*���� 9O����ʽ�'��s���z��ܾ�5��<���8��5e���&L��<�&?��#r�F���8"�q'�����G������a��;�1�ǵ��Elǂ���S7	_�k��
tNwc��j��T�������u������C���5��S��լ��ɿ��Iq(�fiVV��j�CR����S3,~�>n��Z���އ�pX��EW�ƑV����+�e��%@.�pZ$ot��F�JF��{;Lo���h���g�z$����ZQ:@}m׃�(�tɾ�Qu��fs���O+�9B@eCe���K4�H�.�?-��{<��
�����H��xX�3�^�ƅ��GR_����'e�.>z��\W#�,��?Uǣ:�s7[ᭌ)�������"�����2da��olG�ݡ�ڱ��"���U�m ѯ$47#E�z�?w9�o�:x=��#�x����)Qg�rY2YQ1Zǚ�+Z߹��\���JI�^.�uW�<��l�1�֚�;ē�����oA���`T���s����8{c�N�u}�D�Up��2��!�>F�ME�?)�יA� .�/��J=��d�ٛ�XI�̗;��Y�d�<���l�#h��f��EXA�[�R�Z`̌��y��xl׸�3�œv8t����'�nMo���2c��Ht13��T��&���{�g�&��:;d?��&����Ŝ��@���$�T˄���������[~�Y�|T/;j�C��HwS�7%�v���6%�"!��S�sS����!��
���2"��W�HZ��?�R�r�����:����sX�&�5@�o��F��>s�t�����g��7�,ƅ�DB#����=o�oKľ�+���]���s2��\�޼#�Zэ#�ߵ�N|��?`ɡ�܌ۦ���x��/���5W��z�L	���~&��z��A�RLͅ_�#
S"�r%�zk����Ȉ��A�����]u����_v+m�մհ^���'�Q�mY;���J�%%���c�v��y��1���B�e���JɗNBh7�83�i��ܚK�n�Q=��Gia�0.��U�Vp����순� �������u�N��՘��7㖩7��w�S�\��2̯�-�"���A���9t�J���s��Y実���Ԇ-@w'kd�ܢ�Ff�1K���9��h��~���1���C�׿?�0^�]zؤ���r����I�Y����:\��syKS:������ʵ�/ݼ��+��P��N�TJ�I���xGȢl�y�ᅏ�Y��R�8� �Gj��g�L�4��-�B������@8����&V�_�&m��\�p��d��k�MdW�
RU#S��䴴�� �E�;P��"������w)��W�j����_�Aܿ�,Sg%
����F�tLPT�vzy%�f�c�Ԇ���d}�+��y�/�&�g*�<&^uV�I4%�&�N�~�#l���,vF�ժ�Ǣ"�NU�$t6<�<@��P^<I��T�3�I@@�h$��=粓�ߖ��K�Z0ǋ�� u7�\A�o�>-�׈�n���a�5`1!A����yXl%��\({K*S�)��������u����FNa0��WV�A�G������� �h?�_��/��(�ci*�����%[��4�f�H��:���\�f�'���_���W>3o����T�©X�&�6�1��$��-�&���r>:�����wt8o��s(�`�Brl�X�T(������r��e�~��!�YvKӦuw�8�kse����3.� �b���w�![��Y4�Q��-JG)b���G֨�8�rP�<�"��C� M�y8���,�q{"�V�����V�XFYG>p��ٱ6eY����4��T>���'��W�ʔ!��y�Oh���o�a�˗<֦������.}iܻ�Ba$a{<���2iJF_���U&|�"~�q���*����]vsJ�N�^�*C:O5��[-��W�ל�+���M^1�/؈p���Z���i.���<Y� یL@��V�&�i1�8(^�k 9��������0n(`��l���E-�zڏz#n��\��������Id5W��ޒ�r�$ ��?o8��H|��oL����j?E�V���B�)���.�<nQd�5	�_)
�Ix�ѧ7�!��=|~�W�!he�l�[���P~Z:�׃��|���xM�5�9����T�����fS�ǭݭ���va�p�Εx�"�Ń�	M�f�:����I4�����(��Vo�I�!�"�f��hb���£kn�~��N�<-�ɥ��&Y�9ו4v�F�$�X'hu�2�x}2��.�����}<��i�4U]�̊a�.�+e�W��w9��K�<���k h1��c	V~��O�$8���������v��)�y��a�mrF>�^]�N,)�°����XK(>�(�[��ק+�~йea����
�@��`� ȇ�f��gh�� K��d`M�&q���~��z�#Ӂ��|֧��3��z��Q5<Pr��"��J�*x�>Z�0����8B�\����ҵ�D����d�m�qJ��ɹ��05!WOU�%�1�q�A�ۢe�X�c��&��Ar(FIen��^����3Γ�ُY�-9C��!�;��t���MuqY]C[�$�5p�Ƙ������R�sp(I�g|��Q���Z�H1�lZ��{�u���@zI��k��q��]/�.Y���MC!@q%a�.Qr8�_�ؿ,�=��7�4���z%��
�����-{��B^E�H����C�-��WW�ϡ�#J�T]�q�X�u�8Ȯ[K�(Mǹ`�'Uwy��6'CD�d��>}a�rcKG�Yؕ�{nӾ^i��qtq�z�z�5�j�6���^M� �*��z�s������u��rv}kE�A�>�cm�.V�D�׼2�5\d�C�D[����[��C^�+�_.A�b�D��/�
�U��H��ͦ��>��UL����.�z��pV:&`����H	9<��bO�EðU��3���>
�*xg���b�N�

xӶ�y�=���^�k6�7�a��7W��b�:Xi�q��/��>]������;D�7��,�U����SK4�~��b��?�,��"�||{h�A��-�k���{�ʨ�kjz�V���P=�B6u�`���|c���Ҝ�n��wDN��h�%�I(q���\�(E>�w�Х�� MD����v���G�����;�is�dVwv�X��K@���=�%Ԋ5�t�g�]-貀;�[�8`��~���V�-L�uO��į��xe�)���r�JHOZh�$��gv�r�m���Bpr6�qwe���2����!unM�C�F6qe��KS�w��]]^%9�	�!����ٳ�,�Q�t�4�@b.5E�6���?
�����=���~����-8I� 0b�v���,��XJ.1��>�A.?�ϦV52�|�u��D�#����h��;�jÖ?<��d�li�~;�=���K"q[/���H"xÖ#��=ۢ�H��C�A���+DK�]E9߽%��kO��g�d=��X�}q�5.Dj��&_���z!��|z}�����_�Lp�Z�m���� J�8wG�XC�˾�Ú��hDM�����n�ю�b0(X�w],��=���"��E�-��FEx����U�t���7j�0�UL1L�s�o�l�e���WʛH��;�]��l������{�{�>T,zL�J�H�v��ﻣ�sb �Qp�7��!���,٧p��j�/�C��*�'�b؞R�wGH|��oh�-�M��xC: �zxE2�e\+N�u��l�+W��-�?T�$AB"%}=�>�-��I!&���8��A:v�A��e�;�����2��� ��Oz�£l/�>�ZA����Ff2���@3'�d$��t��d�Mn=		r����57�i� ���R٢�~�u����s�G�������\N��T|nJ��)(�o�h��kB��ډ�s!L��HB� �E��T8J���t{P����_9��l����%j,?u�W+W�Ȩ��qm����#
�X���`	��:J��6��c�]��8�%ļ��F|mk�uV�R${��vT��9��YA�fC��X�m{Z`J�{�Ϗf*(��bN����i�A��~�Li��Dk{\���V�N]o|�[y2Iٟ�zΟ��ۄ�We��M��k�� ��^d�%z��� A���x?eG���s�%�wD�m����Z*�\�O�����Lv�d�R����=��X��w�n��]�>�~���d��WE]<]΋���]uO~�j1��v��G��K���9���gT<ms��JC�n����3X��%Yo���S�+��{��D ��Gߝ��;g2�B���Մ�N�0?Ov&�����W]GnӁ[f�y;��pK��on����P�pD�<�ٸ>[kg3/�q"��q��=h�"i��᷅|g��p]LB���`8��yW%���c��7�_��R�S����h��Ա�q|Ȧ\
�[=4�����]�;��H~�x0�EW=4��O��P�s|���\rY���4��� �����<%Ar]_�_��~�$<B�6'�y�d̎�� �߆<�m& ^N�������SOD#�E���K{s��G�[Xeǋ���;���F��'z�#m��������#��H.@>���h�7��V~r_$8�n̦]����j2�b���i��:���$\����#�M�1;椽p�q�5L������T�o�N������)^��%�i�;Q�7n�w�4޾�N�go4�Qt$X"�0Yq$P<JQ�7a���o���㈧�)�3�j�u����cH���7F�@�nI.�*�ժ32�-�W�N��T�*�$����4j������$�r�y����F�Ѩ��Ú-G��d�fÝf�k�n@9ƞ.!��a��:���q���(ĵ�/ߏ��i5<�wL�Q $���$;��<�J'����W�05�zÛ��0-��R��x�=W���^̂����LC<=�<���o�|�l�q"}y1e�\�}�F���[5�u[��K5�H����B{Ƿ���Ś�=洩�ȇ�Z	��?�����S�u��{�c�z�Si_ɝ7�����Ajl̥!_v86y��̋��]J��J�FMzsH����-t�㔫��-�q,�A����l>I��%gw�B�D÷�zk��:؏/�c��vDY�<Wb��Ee_��.�º�ޘ���5n/և�}$L�嫻���E\`���Xv#��C��������|��@�Ԭ���ײG$�3km�JMDD��B����=R���VCaЫi�nSA����6��mb�9�Q̭������@�йV�ZFff<���ݤN�Ht��`���3���|5cA��ô*L �[�`�����R/噸�t�,���4���X�7�T�����F'���,���5u�2Xli�kM̀Si��O<���͛�i'+{��#�~#�Z{�N�[1���|��$�pيtcn���,хbN�����Ѵ*�z�Z��-�ֲs�էit�}o�[WS[�lO�5`B�~�^R0G-ח�Pl7��j���/�>�c���6�+�G�\�&U�դe�Hr�5�i����iܛ5���7^��2�^�þ�}��IB���Q�� -�S$t7�sm<^j����ЯwUpŠ���G[�&�j�uE�]�$j���Z�����.b���<��[ROU��g��nwѫ�T\�v�,8XK�q�G������ؒ��QR��R0\/�w%1�C�n�y.���l!D�l?4�2�b0ADq	b�,8Yu���Y"�k��Z>K{i)�?�7b糂�g���k&�O��')��wm*�\���4 �{��/l����1��h�|�]�|9b_�v����>캜�����'�y�BO��nc��\��аX�?�]���U�ׇ�������`��ŋ��� ���������{"�2n��G��}��.6��r)AΜ���6s�Kͼ��u?L0P##�����QT�x�DC�}�q�;w:ڵ�"3�x�u�ͯ�
�S����6����y;��	�[Y������ٿ��5up��O�DQK ��x�A�[a������������_��ZN�D���|nꮶ�{)�����wX��P�w��X��r;< �t����4�v��`8+�M��""�O-�]����=��I���d�*f�"������0zo??aaFTﲝH�,�i 銂7`�QtUֽ��ޓ�BѪ�����p�%�/���);�}:����jb�;B#Kx3
�[��	��_����������g�'�lҭ��R����=N@�;18Z���V$�[������[�.Ì�Wb�1M��������ɩ�~QȊD���	RE�����ɽe:4Br(��^�V���6����(G�0f�[�-Q8�3C��(I\���D�[�P�=6�������t9r&9��09��%;WP)+F����NV�=��^(��ȵW�:�U��/�*��J>}˴��W+�|,Z z��x/έݱ��NR�Ur+�T�� �Ƃ,����k���~"k�?%�V�,�[�Վ�]*C��s�ZV��q���o{"�<y�m'�����՚��;�S�v����Z�\/w���_Ʋ�,�9�^7��_�UQ��]!�X"l�Es8���a_��O9����*��;�\�s�;�@�x� l|d.%������z5pp��u�6c�^<�m�H��d V]�_5��G~|�pOzN��S�="��֊eڻ��o�}d�Y�q�u�M4Gì`P�W��<In�3Ja��IN�J�d։7C�M4�&c74���M���K�h"�="��m�L"��z� So�܍�yd�:����v�fV�q�
s�x���ьT�y���]� ��Ӽ1g���y�#;e��(����������s��7�y���>���������o��r���V/�Py�ޛ@�	�p�ת�7����^ȳ{�E?H�)��/�!q��t��*u��m`T� ��T��;�"���qn�W��_	8�b-�����NC+l���zݜ�@�.I�8�o8qc���H�$���>����u�;�1�W.\oz��tq��;T�PR���2)�3:���8�	;�v�s,�d���ob��A?��C���6@`k���������a���z(�z�Fi�;ء������;�ߛ^2Y�Y�0��!�nq��S��x�5yWC�0gY5t�k�)M�ݗ/g����4�6��hg�d�Gt����xd������ξ	�������砒Qj�@���ϓ�Y�j�4�Sƿ�E�{�6�61̡�ڸ�̮������\��Bx���!��f�Z�Q�*z��#T��BP��@!9�1�tPp�Lf�Ha�KNy��lX������{� �N�GSL#!�"$U��ը�mE>�'Wj�o�
���Q�V�8*e�=h��E��q���UZǤ�VdEX�i�)�.�jTK!��^�[�%���$/�؜��>�����j�-ռZ9��Y�� h��\��V�2C�2�1��nI��F��k`�m�~X(������/��)��Jӗ;I�fߒ�x��k�W�W#k��R&_�l�u0���c�c5�^"��'�����eH�B�����[���V�F5��_7TnV+��ؒ���粢��#��82��ε���mQq�q�{��}bؾ 3�"b�ri��E����RR�Rx~[�sྩ� '��@��A������vK��ˆ�0R1���9}��ш��J��dݓV�8%}���ŝ�>��4�Z�VHR�����DAG�o�]�ļ�#:����i��:ج��	��!�ʹ0�~���A60C�SJ�"�"�v�J�T&)*[�&�$�	W��'aߵ.�kk%�7��r���K���j�G�<�HŶ���N��?�ԍ2�B���e��]}�,`�2d�iC�8��� 7���ҥ�e�1#q��=z�9r� ڈ���r�_Lh�ڶ�Z[~@����3LϲZ�
���]P4QyU���<2&J���T��CMk&@��F�zq��~F�d}_N��~����1g����6a�!;��%�g"���kb� ���{Dn�o%������>������ ��iT#����(vƃ�f9^P/&[���B�o��?c�fd���z���&Պ=�w3h���H�"��k6x4��Wش�x����z�>T��~l����'�ݓ'�K&?c�@y��ʮ�q{�7���ԑ6~��>ͥ}��8�+�?a�"�~9_d�O2�<��D�{j�@6]|�6�1��H?�P�f7ׁ�:à�C��r:�lIBuۺ-E;;�I�.\�����ce�|ȫ��gA*���/�^�Y���bi{��x�h7�*�mk@`+e�9�1��-'�"�,Qם�+Fo��X	e�,Q�L�u��6�G��88=�����r��B	�T���7��6�.gb8@�L}����^VR0AP@�W�&��&����WU<vKu�Q���luY�{ 7xi�ាy<<jn��E3^��J��a0��0��w,��n�ܷ^.�\�$�	�. 5�E S�8�nI	`��������߷o�#��h�5F5���W�\B�{��;I�o����U�qO�Y4�� ���o�-~�u�.�M���*I35!�y�W���Z���)�ȇ��"�c����FMm��#�a�4�{r�|�	���-�\��ʑ��?����Y������^P|-ʗv�3�Y�q~ױw��� �4�-Y��vd�Z��CƠ�Jc���eP�ԥ�g��!��K���M�k^L�NǮO �f���u��>M����*Sa�(c���d�r��d;���� \�G�!����U�2��V_ĺJpRH�[)�@�j��,���2�3��u�{`����^���{҈%���ǓN�+�'�RT��:�"� �g�ab�5��=�S���>u���Fe�Z˟t(��������1 ����U�S��������O�iBL��pm"�ʡh*�F"��9���>kɈ|t�h{%2����+X2��s��@�yl��u%�2�,���P�ٯ�� Zo^�d�)�; O��q,!t�B��8��z�b5�$�����Xm|�$�������n�W9�B� �_iƯ��|��'��4�)0�C�Y(�6:|q`���w!9�(�(%|{��^_Ҋ6k95C}�䥉{�r��s�xu/�^(�:�|�����*P����� ᑽ�mۀťD5/0�*����WӦ8l�ɳJ�}q��K�B���s9�,z/W+|�:\%+�B��+mS�ڶ$F@C�P�!;�2r`�!e P�;b�eY�t1��Ȉ|�ۢ���No۲�|�Ly����B���`���z�b��S3,���  ���Џ�p|�|OY�
H��.����i��ΥI<���sU-8��w�"��E�z9���j�������I!�.Lk3(�c�%4�����{�o����ŀu�d%[m��n�!�ytƍ �4S�S�I�Jth���&m;hO&�^\k,G��wX	�����M4X�ݼ���_�z���C�{�vh������*��(n�d���5^�{ci����\Ԛo=]AD� &+ҥb�@�kD��S-ej�C�c@��<$��yw��i�vڷbC6W���@:q!=jC��n�~�zT}�Z��������l/`�N�F��V|�07C�V|B
=J��{��'06�q^*��W�/ ��xm������P������ؿ#��QH������d;y���7��O����Z��Yƃ�^UH��O6��f��Ej���������t�ن�R$E:;����׶��t񡺮D9�ׯ�i9��!N9JQߑ��� ����W��6}�țh��d܅	dl���F�ҧ�y`l��c�M˯��/S|B�ò,�0`�����������BC`:a볞�|��/8?0�z�\��N�u��� ��ͪVD:a�3�LN���d��������IĠ�f⥥���'렂�W�u5�=m�P@�  ]���D����@(Ҥ��	�(�MZ)1 �H���	�!�")�_ ���|3w�G�y���}�{2ss����-�C�]W}JlV.��]��N�s�N��<�� =���AZM�G�Y��=��n����5��;�x�t	M�N'炌�=������|,�3��5@����E�kfM1{p�dZ+b5<}\9�|���эF: `s�c��ﷵx��\�>�X0h�;�o"��S֡������=X��#4.�2=�p4!�Y&�+G��>Q髡×>�.	<.�X�ᛊ똒wx��eB}9��SBߐ�E�ޙsy:o�'C�=���}�T���5��Z�����X��-�-�n�=�`ü��笯����M�ި���e��Й�Wf��7!�+н��� ���ܚ`�arf�(����?�C?Cẝ�~4�=���H^{!�0�LR䃢XG�oj�����L��E/SFo �?g�f�Ǉ�}�z.�e��QR}c��9��o��i�T4ʎ����� 2�^}�>�CR�)h�f�Q�w��o#B񷎚?ub^���k����
�x�U90��q�>���`�z�1p���r�������&�Q�2�o��RKX�Ӷ�)�����ix�.�]����M�g�w5��V�eR�̎����(z��eS��~�X��ؙ��;P�]���h@��u]�(t����d�=�G�r{�)����}E�^񣓐O�Y.4n(;+�>�ѹ5=��R`F���hµ`/� *H�&uC���p��s�m|B�-��$��d��9�]Q����SѠd	���o�E������are=6���Lwf��w�v���C�Ks�|r����-�����Q�������z���@�@��"c������[�8K�[f�
��W4~V"L��6����k�M��yB�'/�wѮ�p��"N�	��?}:�������h-]1T�-�k��U4;I=� o�^�c�+}�f����y>�2b����s_��qe]nO�i���ޅ��>h�����>��J�1ǡGXXp|1a��H@��?Nr&n�>��&������0_�W^��d<ώ�,���s;���55C��yi�A����'�����ZEt�M��Xr�3�:�/��w!�U�T��1XD2�H��Z|7)ѿ%+y;�X�zFE�t@��S��h�1٤�1�X�-�3�u}"�O�nm-��2ڏ<��՞a�@W9��x��&��=}��G&K��N/�E"}F,H�k��Z�X����aNi���=�K�U� F�/��ך����a�z�R���W}C�[\�)�����v��ģŻ]>�ˈ ���{e
�lM�~7n[Y�\jm����S��ipv*�;-�� ����R�wz���V�x��fۿG�4�*�U�	Ov$�����A;�A��ϝU��#
ő�RU����A˓����[>��	������'�c���]nQ��g�'�ߊ�\�6�Ӟ�ү���1���W�:2���$4mk��sEM�6X����h��h��r� F?���T�4����*��{����[3�u�6֯�cM�x��8�,hp�LÕ?hm'�q�/�?7�:�ġQ()cbP��f�-н:�t�h��I7��%��m�����9��k)��$��nH�%�f¦_$���1!�֭��U^����
\�*�X3 b!�K,(�}ӨM��`�ű��Z����J�ݔ�@C�5�׷ǍS��w^A�������G]��q���ߐ�Ai�������ܙ�[�$��4[���;&�(@jʥ�2��U�5�{BB��r<g��Z�%�[hX���6�[�R������ɏ���l���T�e3h��m�<��n{Q�m�F��:J��CצcGۼ^]��c����}z��]����{�8��Q�1��
���u֫����ϧ�I��=�_ZX�o�mճ!�ku7n�,���)
v��\�X�� X��I��ۦ4���aX+s�Rf�g��%���؈��%�������`_
0�^�MP���7�"{����}�/��_��e`P�k����}L�� ѱ�JպSrȒ�h�{D��R����ɾ^��\��u�r�CZ�R/$v�,�i��z�u�/ﶒw��\�(�V/L��T���~�T�$Aw{��q�,�T�N=F��^��<�ɍZ�t[�w{9���*5���o'�zԮ��V%���ID�%��@I
@��ݹ�=�Fl��h?��� m|�{Cͨ���[��V���#<�z������$��;P�<�����[H��<Y�;Iا?i��~՗8[_�p�Wj%����ތ�B�ϻ�����T�T-_�.~�8���F�N�}F�]dz%fH�O�~�*\V��ݰDk�c�e
�-�����D��3��y�[u,ٳ}�j�ЦXY͌��gBC㈏�b �ہ� *�!��(��d��s�30L��+/���^��A�yu����� 9�։\mf��Vm��f(��Ob�Wr���1�1�1��0�u8� V!ީÕ~s��ukz���,}���MO�X0�?J^:f���.'�`^_�ݧ8֡4�]]e#�rj�:���
��45,���R}`l�J�x���_K�I��6~Sq��"�9��8�0$ S�aC;�(b#����{��P�]0�}�al�U��D3_����i���!�N�Qխ��AY��7�+�d=N���Hn#�a׺��~�$�ݶ���a�t+�G;�8vr=f�ڑ&>ji�/�L�ߕ�h=в;��2F�k��<φ2LB��Օ>�"�4�2T�U��ʀm*՛u���O�Ǥ��)��X)��G����˺,Y�m�ų�;S�S���1�S.IF�@�����ݵ�{t1pՏp�0*/����p�C���K��!��]g�}�PT7�͌��w����yH"X�;���$G8m<}�͋&>�aj�.�H�������~{��~��˙�U��R_�s't�^�ݣ;iyOƋ�/ �O�S�6�;�H�uc�˝L~��Ā`�:���|������o��\"�4�ީ	�i�{_��8�0��FA!�&��
P�e�ؽ�ڦl��#���pVd �gY��7�ezoªJe�ƅ��E��ƢH�'1R��}[�\`�NMz�+��3�>��pЈ�_g�h:�����=Q$�v��
Z������(�>dh�;In�Y�Xe���{�@��=H�~��z��V�*9��#}���|o��M����MFs��ӂ/f�-h���i}�^�L���g���CK/��|@nF���Z'l�0��^B�-�{P�-�]4Ƕ�,IG�_��.�t!�i1yVY�q����^�ڧUi'��
v��K �25_U�1,;�a���9v��f@~t���l����^5�ӄ����R%�+�x����E��ڎ[y�2l�N�1Y�f �Xdz�f���~^fNɲ�Ӎ��\t���)c�zP��r��~*�6Y���M�h�?Q�H��lj�p��"9��1!A�,)���}a�>Sm�Q[�Y�C���$�|6�6Gy� i`��DT�nO��|�:&c��W��"�8�0��F��U�����k!����wV�=*�^�&4q/P��'u��v�%�-2��!�3�W��7�r��i�Y�o�|�d�p����ٛ�PD��{5]�e"��广�`����� �~W�k���ϣ�����4�nW�zw�L��f�J~GM�~A�r��\�\f�S��c��"�� F��=ψm����+J��@���!
C`u�<�6�!�:E3N6^0�2�1��*�ˋV)O��j>"��*�ן����`��/�;�
��3��8��
Ms�nltY���<T�?/���������/���<��0]L�|�M{�E�"�y��3ղ��f�Z��aԾz�_v�Pq�_Xxq��Z�aH0�y����Q#$SC��E�^c��F�G����\�����R�7 �
>���0c��UN���5��k5�؛e���ɨ������7����`l�M�M
���g�/c�)l����9�	6:�4V.�����zDl��:+��o�r=�܁<�����`9*Kt7t|4:w�=�KE>-�i����J�>θ�cB�@�!��cz��0G��RTeu��u^�C`k���>��%SM+�N񣴹IQ��l=\������`n�6#T�V�c �y7�R�%�9�r�&K�6�A���,�����k5�Z�M��L��!�;a���v���Z�Q�%���
Z<�@�2�zS5��N��@Q������m�RU2��YOb*���0�[�2i�6�֬ }a>@K��i���M���[0��C,�1�� P@0�h�EK��~��ˋ���/��f���Q(��Ԫ ��2�$�[0�M+\�M�+)�T/_���,�`���%��v?�W2m--*��M�~.콸٢�ww���=��SH˳1���dԢ���K|T7HrO ��^�)�fY�D)'�P%�$ٖ���P����V�*+�FF�g��E�Y�T�T�P�|�*�n���=�S!q����g3�����ܢ��T��/sl���2��9l��2�٩�-�e���;�
l�iA������G.5���&�Y^�r��E)q��e١Xo��b/]��'�F�pK_���;����oh�`��HjƎS�5+<��U��d����}����YB9~JDin`=�Ǘ��שϽ�h(�@�Z�U�u�<_�C/��r��q�?��L��;J�mT�&��@�^����~`*Y�K��CPF��H#�r};+۬��v��ճ:t@I�QW;���p��gfH�Et���D^�F}�^䜒��77齩�~΃؊j���\4�4]
}47I�gc���֧7�=5c�ɻ�VJ];8�EU�_;Oq--�=/�Y����?R5�7hp�ܺ�\�]	�Q�����_FM]�W��&�h����`�b+)e�蔟"�`��C3%�7����"L���QQ�vk��;|��!�j�Q]�pn1ع�*�m`�H�ʵR�1�Q-*�]���o�4-~�siEq��IZ�w��&2���6x>�غ�х(V[?�c��H]��X�U��Q@��d
�����)�L�U�����?71\�\X3;s����]M%w��mi�~o6Sr�
�G��~X����+ &k�k53E����>�F�k)@�~��`��-1�'hK�R�t�o�������j�J'��h�bG]�*d.e@�;HM�z�z�M6�I������ے�����`������
_�\�TB�QlG2�?�ɹ��U��$����>�������M*S=�0oۚ~� �%8h��̒�PpT_�堣���o��Q��(���q���\�4���
��vVHǹK�&�
�]�>c����>!��ݘ�'F�J�s����-�Z�Ws-��ju=W����X��Ӷ[$M߂%���?�`�濾�5�@s�
����!��r���0#�B�e��@Z�z�r˸����R*o؜��j�n�ZsI�1L���ڡT�H�����403��l��\p����)���OȨ�˕��ڮ7�S2�^�V�U+^/�p�ȉ ��愊k�A�ߴ�y���$�A�A���L�����	a1�G��#�Ob��~c5�~�_�n�Z@Y��i<b�H�P�d�-U �:pi��E��;nU�Lm���КGn.�^��K�UAmt:� `��մ��9�?�Y��<ψF���_����� ���C��Ԭ��PK   w~�XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   x~�X�I��J  J/     jsons/user_defined.json�Y�n�8}Ëv��H�'I��I��� �H*�H�,5�}�}�}����؎>B�f1X���X4y�%y�!�Տq�}��G�r��[��$uv<u�*�R�O�@˪������?<=��j�,�e�f�O������e�w�8���<3YZ��b���ͤ6t��s���M�	|Sf#�1CR�$�iL#�"-RH��Ə�2y�,'7헉��S����"nI���I�g8F��2��q�B�������L3�a��gi���~����$Y-��q�XU��S]6�W�c�N���*�i���3;/���rV�UR9�!Y@aO�~HV���g9y	K�Б�z}:�4?=��tÒ6,�]/������^Xچ^�Wn�^Xֆ�`ٔ]���6��B������0�~޿YA4��Ae�b/�kh�UmP�:ý�a��/1I��iE��F�Aۤ�~�?c��mJQ�؟�~�6��_��D?h�Oa�'�
:?~ߏ��(�	{2����	 iӊP?�!��6��=!���ᾰ�D������'-�8�_�~}�����Q;�,剪�Q��U�U���9F�'jЏڦX}�����8��'j� Ҏ��{��Ӌv]���]���
<Q���:/�
ܺ������1���F�U��`��\1��q�b1��=����2�/��<[��H֩�:�X5����!�i�v�EYg�%������}�x�g�g��\�:Y%��=���KY�[_���鳨�2֦(sHL�L7����540$K]Z\?�SV�A߹��IM򲀯�[�ͽ��s7�� �"��U�`��).xD�fa�,�`��b( �֜ɀ��7�
��9'#�mi�r�C�E��&�el�v{'k��S�uҳ�yRT���C�UW���7R6�e��V�����6+�Eb>��l�lR�mg+{��ٿgC[-kK��Q����"Y?� ��?����y!�A[.lLG�|�˳2��pf����w��oN]�Kmv&E���V���?�zgi1O~w[��? ���qV��G��qș�m-�QX�)r1�4��At;����	�c����<�:�ˤ]�?=}�����ك��|D�l��6� �ӰA��(��)�8%"�h��8D�RA%qVך��y����0D8W��!e`)�@Z��A'�w+%�M�9�o�%޿f����	�2 B���ɇ����`�2�k#X�#������o{TDc�++'Ƿ��}S$�qu:?��G�EV&�Pq��=�.����XԾ̆��[�>;ߣCpeA���:�쾌��{��O�S=i�Yj�j��&����.`�� ł���ETs��Ș	�b!�ۉ�e���ʢ��2=_��s\��2���!r�p䨍�!�+�XQe��L�8�T(PhX��0��S��Z�=d�O%��S�Ŕ����E��`Ji ń����k%nhT��Em@�6U���r8�x�:��ma��g
�-%���#�0�?Cj��+ӷV�8�\!��*a]#J�#�q�BƵ;��AjpP��V�+�JVE�wVlj�Kj�"@���	�Z�K,�\e��%���&�(�Q��VEpB&���A�5��u�Ж�J�U���r'h�xZg���]j_t���� �����}ݾ���'/X�Кd-��Nk�{շ��ՆM���l�E(��E����h��e�	F&�J�wU�
Od5ϛ-NZp�f�����l��]�c�<du�UN���MxJ��S��V�G�K����9/"��.�ѯ:���Ob�!��I�ekG3��C�U�k�Q�G�-@�%�RE8(�A�pP��"��[E8��=��^�������PK
   x~�X�c�-)  Ǆ                  cirkitFile.jsonPK
   w~�X����7  �  /             Z)  images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   w~�X��Q"�  �  /             �:  images/6e6351c6-f51b-4efc-b2a4-a37f35def552.pngPK
   x~�X�x�LA �h /             �V  images/7f6d2589-4c6d-4619-9f3b-04025fafdd34.pngPK
   x~�Xd��  �   /             � images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   w~�X�&�}[  y`  /             )� images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   x~�X	��#u } /             � images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   w~�X$7h�!  �!  /             c� images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   x~�X0%�a�  �  /             �� images/d63f6a48-eabb-43c6-9b21-e1ae45e934ae.pngPK
   x~�X�tԿI� � /             �� images/d8a77cc3-1409-488f-923b-bd8c8826a526.pngPK
   w~�XP��/�  ǽ  /             � images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   x~�X�I��J  J/               ic jsons/user_defined.jsonPK      $  �j   